library verilog;
use verilog.vl_types.all;
entity acc_cosim_wrapper is
    port(
        \_RESET\        : in     vl_logic
    );
end acc_cosim_wrapper;

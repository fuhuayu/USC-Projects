library verilog;
use verilog.vl_types.all;
entity acc_csp_gold_sv_unit is
end acc_csp_gold_sv_unit;

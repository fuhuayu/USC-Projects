library verilog;
use verilog.vl_types.all;
entity middle_finder_tb is
end middle_finder_tb;

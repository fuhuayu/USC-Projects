
module TCAM ( reset, clk, DIN, EN, WE, match, match_addr );
  input [15:0] DIN;
  output [2:0] match_addr;
  input reset, clk, EN, WE;
  output match;
  wire   n84, n85, n86, n2999, n3000, n3001, n3002, j_3_, n87, n88, n89, m,
         n250, n251, n252, n868, n870, n873, n874, n876, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n895, n897, n900, n901, n902, n903, n904, n905, n906, n908,
         n909, n910, n911, n912, n914, n915, n916, n917, n919, n921, n923,
         n925, n926, n928, n929, n930, n932, n936, n937, n938, n939, n940,
         n941, n943, n944, n945, n946, n948, n952, n953, n954, n955, n956,
         n957, n959, n960, n961, n962, n964, n967, n968, n969, n970, n971,
         n972, n974, n975, n976, n977, n979, n983, n984, n985, n986, n987,
         n988, n990, n991, n992, n993, n995, n998, n999, n1000, n1001, n1002,
         n1003, n1005, n1007, n1009, n1010, n1011, n1013, n1014, n1015, n1016,
         n1017, n1018, n1021, n1023, n1025, n1027, n1028, n1030, n1031, n1033,
         n1034, n1036, n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1049, n1051, n1053, n1054, n1055, n1057, n1058, n1064,
         n1065, n1066, n1067, n1069, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1086, n1087,
         n1088, n1090, n1092, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1113, n1115, n1117, n1118, n1119, n1121, n1122, n1128, n1129, n1130,
         n1131, n1133, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1151, n1152, n1154,
         n1156, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1178,
         n1180, n1182, n1183, n1184, n1186, n1187, n1193, n1194, n1195, n1196,
         n1198, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1219, n1221,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1242, n1244, n1246,
         n1247, n1248, n1250, n1251, n1257, n1258, n1259, n1260, n1262, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1279, n1280, n1281, n1283, n1285, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1317, n1319, n1321, n1323,
         n1325, n1327, n1329, n1331, n1334, n1335, n1336, n1337, n1338, n1339,
         n1342, n1345, n1348, n1350, n1352, n1354, n1356, n1358, n1360, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1395, n1396, n1398, n1400, n1402, n1403, n1404, n1405, n1406, n1407,
         n1409, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1441, n1442, n1444, n1446, n1448, n1449, n1450, n1451, n1452, n1453,
         n1455, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1485, n1486,
         n1487, n1488, n1490, n1492, n1494, n1495, n1496, n1497, n1498, n1499,
         n1501, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1512, n1513,
         n1514, n1515, n1517, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1531, n1533, n1534, n1535, n1538, n1540, n1542,
         n1545, n1547, n1548, n1550, n1553, n1554, n1556, n1557, n1558, n1559,
         n1560, n1561, n1565, n1567, n1569, n1572, n1574, n1575, n1577, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1588, n1590, n1593,
         n1595, n1596, n1598, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1609, n1611, n1614, n1616, n1617, n1619, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1631, n1633, n1636, n1638,
         n1639, n1641, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1652, n1654, n1657, n1659, n1660, n1662, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1673, n1675, n1678, n1680, n1681, n1683,
         n1685, n1686, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1708, n1716, n1781,
         n1844, n1890, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n238, n236, n235, n233, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
  wire   [23:0] rank;
  wire   [127:0] mem;
  wire   [23:0] matchN;
  wire   [2:0] last;

  DFFSR rank_reg_0__0_ ( .D(n2073), .CLK(clk), .R(n2786), .S(1'b1), .Q(rank[0]) );
  DFFSR rank_reg_0__1_ ( .D(n2071), .CLK(clk), .R(n2779), .S(1'b1), .Q(rank[1]) );
  DFFSR rank_reg_0__2_ ( .D(n2070), .CLK(clk), .R(n2779), .S(1'b1), .Q(rank[2]) );
  DFFPOSX1 last_reg_0_ ( .D(n1899), .CLK(clk), .Q(last[0]) );
  DFFSR matchN_reg_0__2_ ( .D(n2031), .CLK(clk), .R(n2779), .S(1'b1), .Q(
        matchN[2]) );
  DFFSR matchN_reg_0__1_ ( .D(n2032), .CLK(clk), .R(n2779), .S(1'b1), .Q(
        matchN[1]) );
  DFFSR matchN_reg_0__0_ ( .D(n2033), .CLK(clk), .R(n2779), .S(1'b1), .Q(
        matchN[0]) );
  DFFSR mem_reg_0__15_ ( .D(n2034), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[15]) );
  DFFSR mem_reg_0__14_ ( .D(n2035), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[14]) );
  DFFSR mem_reg_0__13_ ( .D(n2036), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[13]) );
  DFFSR mem_reg_0__12_ ( .D(n2037), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[12]) );
  DFFSR mem_reg_0__11_ ( .D(n2038), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[11]) );
  DFFSR mem_reg_0__10_ ( .D(n2039), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[10]) );
  DFFSR mem_reg_0__9_ ( .D(n2040), .CLK(clk), .R(n2779), .S(1'b1), .Q(mem[9])
         );
  DFFSR mem_reg_0__8_ ( .D(n2041), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[8])
         );
  DFFSR mem_reg_0__7_ ( .D(n2042), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[7])
         );
  DFFSR mem_reg_0__6_ ( .D(n2043), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[6])
         );
  DFFSR mem_reg_0__5_ ( .D(n2044), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[5])
         );
  DFFSR mem_reg_0__4_ ( .D(n2045), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[4])
         );
  DFFSR mem_reg_0__3_ ( .D(n2046), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[3])
         );
  DFFSR mem_reg_0__2_ ( .D(n2047), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[2])
         );
  DFFSR mem_reg_0__1_ ( .D(n2048), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[1])
         );
  DFFSR mem_reg_0__0_ ( .D(n2049), .CLK(clk), .R(n2780), .S(1'b1), .Q(mem[0])
         );
  DFFPOSX1 j_reg_0_ ( .D(n1892), .CLK(clk), .Q(n84) );
  DFFSR rank_reg_6__2_ ( .D(n2052), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[20]) );
  DFFSR rank_reg_6__0_ ( .D(n2054), .CLK(clk), .R(n2780), .S(1'b1), .Q(
        rank[18]) );
  DFFSR rank_reg_6__1_ ( .D(n2053), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[19]) );
  DFFPOSX1 last_reg_2_ ( .D(n1897), .CLK(clk), .Q(last[2]) );
  DFFSR matchN_reg_7__2_ ( .D(n1894), .CLK(clk), .R(n2780), .S(1'b1), .Q(
        matchN[23]) );
  DFFSR matchN_reg_7__1_ ( .D(n1895), .CLK(clk), .R(n2780), .S(1'b1), .Q(
        matchN[22]) );
  DFFSR matchN_reg_7__0_ ( .D(n1896), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        matchN[21]) );
  DFFSR mem_reg_7__15_ ( .D(n1901), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[127]) );
  DFFSR mem_reg_7__14_ ( .D(n1902), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[126]) );
  DFFSR mem_reg_7__13_ ( .D(n1903), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[125]) );
  DFFSR mem_reg_7__12_ ( .D(n1904), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[124]) );
  DFFSR mem_reg_7__11_ ( .D(n1905), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[123]) );
  DFFSR mem_reg_7__10_ ( .D(n1906), .CLK(clk), .R(n2781), .S(1'b1), .Q(
        mem[122]) );
  DFFSR mem_reg_7__9_ ( .D(n1907), .CLK(clk), .R(n2781), .S(1'b1), .Q(mem[121]) );
  DFFSR mem_reg_7__8_ ( .D(n1908), .CLK(clk), .R(n2781), .S(1'b1), .Q(mem[120]) );
  DFFSR mem_reg_7__7_ ( .D(n1909), .CLK(clk), .R(n2781), .S(1'b1), .Q(mem[119]) );
  DFFSR mem_reg_7__6_ ( .D(n1910), .CLK(clk), .R(n2781), .S(1'b1), .Q(mem[118]) );
  DFFSR mem_reg_7__5_ ( .D(n1911), .CLK(clk), .R(n2781), .S(1'b1), .Q(mem[117]) );
  DFFSR mem_reg_7__4_ ( .D(n1912), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[116]) );
  DFFSR mem_reg_7__3_ ( .D(n1913), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[115]) );
  DFFSR mem_reg_7__2_ ( .D(n1914), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[114]) );
  DFFSR mem_reg_7__1_ ( .D(n1915), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[113]) );
  DFFSR mem_reg_7__0_ ( .D(n1916), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[112]) );
  DFFPOSX1 j_reg_2_ ( .D(n1890), .CLK(clk), .Q(n86) );
  DFFSR match_addr_reg_2_ ( .D(n1844), .CLK(clk), .R(n2782), .S(1'b1), .Q(
        n3000) );
  DFFSR rank_reg_5__2_ ( .D(n2055), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[17]) );
  DFFSR rank_reg_5__0_ ( .D(n2057), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[15]) );
  DFFSR rank_reg_5__1_ ( .D(n2056), .CLK(clk), .R(n2782), .S(1'b1), .Q(
        rank[16]) );
  DFFPOSX1 last_reg_1_ ( .D(n1898), .CLK(clk), .Q(last[1]) );
  DFFSR mem_reg_4__0_ ( .D(n1973), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[64])
         );
  DFFSR mem_reg_4__1_ ( .D(n1972), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[65])
         );
  DFFSR mem_reg_4__2_ ( .D(n1971), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[66])
         );
  DFFSR mem_reg_4__3_ ( .D(n1970), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[67])
         );
  DFFSR mem_reg_4__4_ ( .D(n1969), .CLK(clk), .R(n2782), .S(1'b1), .Q(mem[68])
         );
  DFFSR mem_reg_4__5_ ( .D(n1968), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[69])
         );
  DFFSR mem_reg_4__6_ ( .D(n1967), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[70])
         );
  DFFSR mem_reg_4__7_ ( .D(n1966), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[71])
         );
  DFFSR mem_reg_4__8_ ( .D(n1965), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[72])
         );
  DFFSR mem_reg_4__9_ ( .D(n1964), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[73])
         );
  DFFSR mem_reg_4__10_ ( .D(n1963), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[74]) );
  DFFSR mem_reg_4__11_ ( .D(n1962), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[75]) );
  DFFSR mem_reg_4__12_ ( .D(n1961), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[76]) );
  DFFSR mem_reg_4__13_ ( .D(n1960), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[77]) );
  DFFSR mem_reg_4__14_ ( .D(n1959), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[78]) );
  DFFSR mem_reg_4__15_ ( .D(n1958), .CLK(clk), .R(n2783), .S(1'b1), .Q(mem[79]) );
  DFFSR matchN_reg_4__0_ ( .D(n1957), .CLK(clk), .R(n2783), .S(1'b1), .Q(
        matchN[12]) );
  DFFSR matchN_reg_4__1_ ( .D(n1956), .CLK(clk), .R(n2784), .S(1'b1), .Q(
        matchN[13]) );
  DFFSR matchN_reg_4__2_ ( .D(n1955), .CLK(clk), .R(n2784), .S(1'b1), .Q(
        matchN[14]) );
  DFFSR mem_reg_2__0_ ( .D(n2011), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[32])
         );
  DFFSR mem_reg_2__1_ ( .D(n2010), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[33])
         );
  DFFSR mem_reg_2__2_ ( .D(n2009), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[34])
         );
  DFFSR mem_reg_2__3_ ( .D(n2008), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[35])
         );
  DFFSR mem_reg_2__4_ ( .D(n2007), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[36])
         );
  DFFSR mem_reg_2__5_ ( .D(n2006), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[37])
         );
  DFFSR mem_reg_2__6_ ( .D(n2005), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[38])
         );
  DFFSR mem_reg_2__7_ ( .D(n2004), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[39])
         );
  DFFSR mem_reg_2__8_ ( .D(n2003), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[40])
         );
  DFFSR mem_reg_2__9_ ( .D(n2002), .CLK(clk), .R(n2784), .S(1'b1), .Q(mem[41])
         );
  DFFSR mem_reg_2__10_ ( .D(n2001), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[42]) );
  DFFSR mem_reg_2__11_ ( .D(n2000), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[43]) );
  DFFSR mem_reg_2__12_ ( .D(n1999), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[44]) );
  DFFSR mem_reg_2__13_ ( .D(n1998), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[45]) );
  DFFSR mem_reg_2__14_ ( .D(n1997), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[46]) );
  DFFSR mem_reg_2__15_ ( .D(n1996), .CLK(clk), .R(n2785), .S(1'b1), .Q(mem[47]) );
  DFFSR matchN_reg_2__0_ ( .D(n1995), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[6]) );
  DFFSR matchN_reg_2__1_ ( .D(n1994), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[7]) );
  DFFSR matchN_reg_2__2_ ( .D(n1993), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[8]) );
  DFFSR matchN_reg_6__2_ ( .D(n1917), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[20]) );
  DFFSR matchN_reg_6__1_ ( .D(n1918), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[19]) );
  DFFSR matchN_reg_6__0_ ( .D(n1919), .CLK(clk), .R(n2785), .S(1'b1), .Q(
        matchN[18]) );
  DFFSR mem_reg_6__15_ ( .D(n1920), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[111]) );
  DFFSR mem_reg_6__14_ ( .D(n1921), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[110]) );
  DFFSR mem_reg_6__13_ ( .D(n1922), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[109]) );
  DFFSR mem_reg_6__12_ ( .D(n1923), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[108]) );
  DFFSR mem_reg_6__11_ ( .D(n1924), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[107]) );
  DFFSR mem_reg_6__10_ ( .D(n1925), .CLK(clk), .R(n2786), .S(1'b1), .Q(
        mem[106]) );
  DFFSR mem_reg_6__9_ ( .D(n1926), .CLK(clk), .R(n2786), .S(1'b1), .Q(mem[105]) );
  DFFSR mem_reg_6__8_ ( .D(n1927), .CLK(clk), .R(n2786), .S(1'b1), .Q(mem[104]) );
  DFFSR mem_reg_6__7_ ( .D(n1928), .CLK(clk), .R(n2786), .S(1'b1), .Q(mem[103]) );
  DFFSR mem_reg_6__6_ ( .D(n1929), .CLK(clk), .R(n2786), .S(1'b1), .Q(mem[102]) );
  DFFSR mem_reg_6__5_ ( .D(n1930), .CLK(clk), .R(n2786), .S(1'b1), .Q(mem[101]) );
  DFFSR mem_reg_6__4_ ( .D(n1931), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[100]) );
  DFFSR mem_reg_6__3_ ( .D(n1932), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[99])
         );
  DFFSR mem_reg_6__2_ ( .D(n1933), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[98])
         );
  DFFSR mem_reg_6__1_ ( .D(n1934), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[97])
         );
  DFFSR mem_reg_6__0_ ( .D(n1935), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[96])
         );
  DFFSR m_reg ( .D(n1900), .CLK(clk), .R(n2787), .S(1'b1), .Q(m) );
  DFFSR match_reg ( .D(n2556), .CLK(clk), .R(n2787), .S(1'b1), .Q(n2999) );
  DFFSR matchN_reg_5__2_ ( .D(n1936), .CLK(clk), .R(n2787), .S(1'b1), .Q(
        matchN[17]) );
  DFFSR matchN_reg_5__1_ ( .D(n1937), .CLK(clk), .R(n2787), .S(1'b1), .Q(
        matchN[16]) );
  DFFSR matchN_reg_5__0_ ( .D(n1938), .CLK(clk), .R(n2787), .S(1'b1), .Q(
        matchN[15]) );
  DFFSR mem_reg_5__15_ ( .D(n1939), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[95]) );
  DFFSR mem_reg_5__14_ ( .D(n1940), .CLK(clk), .R(n2787), .S(1'b1), .Q(mem[94]) );
  DFFSR mem_reg_5__13_ ( .D(n1941), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[93]) );
  DFFSR mem_reg_5__12_ ( .D(n1942), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[92]) );
  DFFSR mem_reg_5__11_ ( .D(n1943), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[91]) );
  DFFSR mem_reg_5__10_ ( .D(n1944), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[90]) );
  DFFSR mem_reg_5__9_ ( .D(n1945), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[89])
         );
  DFFSR mem_reg_5__8_ ( .D(n1946), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[88])
         );
  DFFSR mem_reg_5__7_ ( .D(n1947), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[87])
         );
  DFFSR mem_reg_5__6_ ( .D(n1948), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[86])
         );
  DFFSR mem_reg_5__5_ ( .D(n1949), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[85])
         );
  DFFSR mem_reg_5__4_ ( .D(n1950), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[84])
         );
  DFFSR mem_reg_5__3_ ( .D(n1951), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[83])
         );
  DFFSR mem_reg_5__2_ ( .D(n1952), .CLK(clk), .R(n2788), .S(1'b1), .Q(mem[82])
         );
  DFFSR mem_reg_5__1_ ( .D(n1953), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[81])
         );
  DFFSR mem_reg_5__0_ ( .D(n1954), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[80])
         );
  DFFSR matchN_reg_3__2_ ( .D(n1974), .CLK(clk), .R(n2789), .S(1'b1), .Q(
        matchN[11]) );
  DFFSR matchN_reg_3__1_ ( .D(n1975), .CLK(clk), .R(n2789), .S(1'b1), .Q(
        matchN[10]) );
  DFFSR matchN_reg_3__0_ ( .D(n1976), .CLK(clk), .R(n2789), .S(1'b1), .Q(
        matchN[9]) );
  DFFSR mem_reg_3__15_ ( .D(n1977), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[63]) );
  DFFSR mem_reg_3__14_ ( .D(n1978), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[62]) );
  DFFSR mem_reg_3__13_ ( .D(n1979), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[61]) );
  DFFSR mem_reg_3__12_ ( .D(n1980), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[60]) );
  DFFSR mem_reg_3__11_ ( .D(n1981), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[59]) );
  DFFSR mem_reg_3__10_ ( .D(n1982), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[58]) );
  DFFSR mem_reg_3__9_ ( .D(n1983), .CLK(clk), .R(n2789), .S(1'b1), .Q(mem[57])
         );
  DFFSR mem_reg_3__8_ ( .D(n1984), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[56])
         );
  DFFSR mem_reg_3__7_ ( .D(n1985), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[55])
         );
  DFFSR mem_reg_3__6_ ( .D(n1986), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[54])
         );
  DFFSR mem_reg_3__5_ ( .D(n1987), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[53])
         );
  DFFSR mem_reg_3__4_ ( .D(n1988), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[52])
         );
  DFFSR mem_reg_3__3_ ( .D(n1989), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[51])
         );
  DFFSR mem_reg_3__2_ ( .D(n1990), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[50])
         );
  DFFSR mem_reg_3__1_ ( .D(n1991), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[49])
         );
  DFFSR mem_reg_3__0_ ( .D(n1992), .CLK(clk), .R(n2790), .S(1'b1), .Q(mem[48])
         );
  DFFSR matchN_reg_1__2_ ( .D(n2012), .CLK(clk), .R(n2790), .S(1'b1), .Q(
        matchN[5]) );
  DFFSR matchN_reg_1__1_ ( .D(n2013), .CLK(clk), .R(n2790), .S(1'b1), .Q(
        matchN[4]) );
  DFFSR matchN_reg_1__0_ ( .D(n2014), .CLK(clk), .R(n2790), .S(1'b1), .Q(
        matchN[3]) );
  DFFSR mem_reg_1__15_ ( .D(n2015), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[31]) );
  DFFSR mem_reg_1__14_ ( .D(n2016), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[30]) );
  DFFSR mem_reg_1__13_ ( .D(n2017), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[29]) );
  DFFSR mem_reg_1__12_ ( .D(n2018), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[28]) );
  DFFSR mem_reg_1__11_ ( .D(n2019), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[27]) );
  DFFSR mem_reg_1__10_ ( .D(n2020), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[26]) );
  DFFSR mem_reg_1__9_ ( .D(n2021), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[25])
         );
  DFFSR mem_reg_1__8_ ( .D(n2022), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[24])
         );
  DFFSR mem_reg_1__7_ ( .D(n2023), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[23])
         );
  DFFSR mem_reg_1__6_ ( .D(n2024), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[22])
         );
  DFFSR mem_reg_1__5_ ( .D(n2025), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[21])
         );
  DFFSR mem_reg_1__4_ ( .D(n2026), .CLK(clk), .R(n2792), .S(1'b1), .Q(mem[20])
         );
  DFFSR mem_reg_1__3_ ( .D(n2027), .CLK(clk), .R(n2791), .S(1'b1), .Q(mem[19])
         );
  DFFSR mem_reg_1__2_ ( .D(n2028), .CLK(clk), .R(n2792), .S(1'b1), .Q(mem[18])
         );
  DFFSR mem_reg_1__1_ ( .D(n2029), .CLK(clk), .R(n2792), .S(1'b1), .Q(mem[17])
         );
  DFFSR mem_reg_1__0_ ( .D(n2030), .CLK(clk), .R(n2792), .S(1'b1), .Q(mem[16])
         );
  DFFPOSX1 j_reg_3_ ( .D(n1893), .CLK(clk), .Q(j_3_) );
  DFFPOSX1 j_reg_1_ ( .D(n2795), .CLK(clk), .Q(n85) );
  DFFSR rank_reg_7__1_ ( .D(n2050), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[22]) );
  DFFSR rank_reg_7__0_ ( .D(n2051), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[21]) );
  DFFSR rank_reg_7__2_ ( .D(n2072), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[23]) );
  DFFSR rank_reg_4__2_ ( .D(n2058), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[14]) );
  DFFSR rank_reg_4__0_ ( .D(n2060), .CLK(clk), .R(n2792), .S(1'b1), .Q(
        rank[12]) );
  DFFSR rank_reg_4__1_ ( .D(n2059), .CLK(clk), .R(n2792), .S(1'b1), .Q(
        rank[13]) );
  DFFSR match_addr_reg_1_ ( .D(n1716), .CLK(clk), .R(n2792), .S(1'b1), .Q(
        n3001) );
  DFFSR rank_reg_2__2_ ( .D(n2064), .CLK(clk), .R(n2792), .S(1'b1), .Q(rank[8]) );
  DFFSR rank_reg_2__0_ ( .D(n2066), .CLK(clk), .R(n2792), .S(1'b1), .Q(rank[6]) );
  DFFSR rank_reg_2__1_ ( .D(n2065), .CLK(clk), .R(1'b1), .S(n2793), .Q(rank[7]) );
  DFFSR rank_reg_3__2_ ( .D(n2061), .CLK(clk), .R(n2792), .S(1'b1), .Q(
        rank[11]) );
  DFFSR rank_reg_3__0_ ( .D(n2063), .CLK(clk), .R(1'b1), .S(n2793), .Q(rank[9]) );
  DFFSR rank_reg_3__1_ ( .D(n2062), .CLK(clk), .R(1'b1), .S(n2793), .Q(
        rank[10]) );
  DFFSR match_addr_reg_0_ ( .D(n1708), .CLK(clk), .R(n2792), .S(1'b1), .Q(
        n3002) );
  DFFSR rank_reg_1__2_ ( .D(n2067), .CLK(clk), .R(n2792), .S(1'b1), .Q(rank[5]) );
  DFFSR rank_reg_1__0_ ( .D(n2069), .CLK(clk), .R(1'b1), .S(n2793), .Q(rank[3]) );
  DFFSR rank_reg_1__1_ ( .D(n2068), .CLK(clk), .R(n2793), .S(1'b1), .Q(rank[4]) );
  OAI21X1 U3 ( .A(n2752), .B(n2871), .C(n2512), .Y(n1708) );
  OAI21X1 U5 ( .A(n2752), .B(n2968), .C(n2481), .Y(n1716) );
  OAI21X1 U9 ( .A(n2752), .B(n2885), .C(n2447), .Y(n1844) );
  OAI21X1 U12 ( .A(n2797), .B(n878), .C(n2388), .Y(n1890) );
  AOI21X1 U16 ( .A(n2666), .B(n85), .C(n2245), .Y(n882) );
  AOI21X1 U17 ( .A(n2253), .B(n2528), .C(n878), .Y(n883) );
  NAND3X1 U18 ( .A(n2597), .B(n2502), .C(n2753), .Y(n884) );
  OAI21X1 U19 ( .A(n2414), .B(n878), .C(n2415), .Y(n1892) );
  AOI21X1 U22 ( .A(n891), .B(n2748), .C(n2798), .Y(n889) );
  OAI21X1 U23 ( .A(n2801), .B(n2276), .C(n2597), .Y(n891) );
  AOI21X1 U24 ( .A(n2812), .B(n2750), .C(n2808), .Y(n895) );
  OAI21X1 U26 ( .A(n2844), .B(n2666), .C(n2434), .Y(n1893) );
  OAI21X1 U29 ( .A(n902), .B(n2730), .C(n2776), .Y(n901) );
  NOR3X1 U30 ( .A(n2667), .B(n2470), .C(n2502), .Y(n902) );
  NAND3X1 U32 ( .A(n2597), .B(n2753), .C(n2528), .Y(n881) );
  NAND3X1 U35 ( .A(n2249), .B(n2266), .C(n2287), .Y(n908) );
  AOI21X1 U36 ( .A(n912), .B(n2878), .C(n2501), .Y(n911) );
  NAND3X1 U37 ( .A(n2252), .B(n916), .C(n917), .Y(n910) );
  AOI22X1 U41 ( .A(n2800), .B(n2309), .C(n2352), .D(n2748), .Y(n921) );
  NAND3X1 U42 ( .A(n916), .B(n2879), .C(n919), .Y(n909) );
  OAI21X1 U43 ( .A(n2929), .B(n2748), .C(n2244), .Y(n919) );
  OAI21X1 U47 ( .A(n2748), .B(n2928), .C(n2306), .Y(n912) );
  NAND3X1 U50 ( .A(n2749), .B(n930), .C(n932), .Y(n892) );
  OAI21X1 U52 ( .A(n2803), .B(n2802), .C(n2928), .Y(n930) );
  AOI21X1 U55 ( .A(n2804), .B(n2713), .C(n936), .Y(n928) );
  OAI21X1 U57 ( .A(n926), .B(n2929), .C(n2165), .Y(n937) );
  NAND3X1 U58 ( .A(n2352), .B(n2270), .C(n2310), .Y(n938) );
  AOI21X1 U60 ( .A(n2728), .B(n2804), .C(n2247), .Y(n923) );
  OAI21X1 U63 ( .A(n2948), .B(n2597), .C(n2243), .Y(n926) );
  NAND3X1 U65 ( .A(n2598), .B(n946), .C(n948), .Y(n886) );
  OAI21X1 U67 ( .A(n2805), .B(n936), .C(n2947), .Y(n946) );
  OAI21X1 U70 ( .A(n2753), .B(n2908), .C(n2499), .Y(n936) );
  OAI21X1 U72 ( .A(n944), .B(n2948), .C(n2164), .Y(n953) );
  NAND3X1 U73 ( .A(n2251), .B(n941), .C(n2728), .Y(n954) );
  OAI21X1 U74 ( .A(n2651), .B(n2753), .C(n2242), .Y(n941) );
  OAI21X1 U78 ( .A(n2907), .B(n2753), .C(n2241), .Y(n944) );
  NAND3X1 U80 ( .A(n2754), .B(n962), .C(n964), .Y(n888) );
  OAI21X1 U82 ( .A(n2807), .B(n2806), .C(n2908), .Y(n962) );
  AOI21X1 U85 ( .A(n2808), .B(n2714), .C(n967), .Y(n952) );
  OAI21X1 U87 ( .A(n960), .B(n2907), .C(n2163), .Y(n968) );
  NAND3X1 U88 ( .A(n2311), .B(n2269), .C(n2651), .Y(n969) );
  AOI21X1 U90 ( .A(n2729), .B(n2808), .C(n2246), .Y(n957) );
  OAI21X1 U93 ( .A(n2955), .B(n2585), .C(n2240), .Y(n960) );
  NAND3X1 U95 ( .A(n2586), .B(n977), .C(n979), .Y(n906) );
  OAI21X1 U97 ( .A(n2809), .B(n967), .C(n2954), .Y(n977) );
  OAI21X1 U100 ( .A(n2750), .B(n2927), .C(n2525), .Y(n967) );
  OAI21X1 U102 ( .A(n975), .B(n2955), .C(n2162), .Y(n984) );
  NAND3X1 U103 ( .A(n2250), .B(n972), .C(n2729), .Y(n985) );
  OAI21X1 U104 ( .A(n2652), .B(n2750), .C(n2239), .Y(n972) );
  OAI21X1 U107 ( .A(n2926), .B(n2750), .C(n2238), .Y(n975) );
  NAND3X1 U109 ( .A(n2751), .B(n993), .C(n995), .Y(n897) );
  OAI21X1 U111 ( .A(n2810), .B(n2811), .C(n2927), .Y(n993) );
  AOI21X1 U114 ( .A(n2715), .B(n2812), .C(n998), .Y(n983) );
  OAI21X1 U116 ( .A(n991), .B(n2926), .C(n2161), .Y(n999) );
  NAND3X1 U117 ( .A(n2471), .B(n2268), .C(n2652), .Y(n1000) );
  AOI21X1 U119 ( .A(n2662), .B(n2812), .C(n1002), .Y(n988) );
  NOR3X1 U120 ( .A(n2537), .B(n2812), .C(n2854), .Y(n1002) );
  OAI21X1 U122 ( .A(n2962), .B(n2591), .C(n2160), .Y(n991) );
  NAND3X1 U123 ( .A(n1003), .B(n2591), .C(n2733), .Y(n1007) );
  NAND3X1 U127 ( .A(n2592), .B(n1010), .C(n1011), .Y(n1005) );
  OAI21X1 U128 ( .A(n998), .B(n2961), .C(n2143), .Y(n1010) );
  AOI22X1 U129 ( .A(n2662), .B(n1014), .C(n2539), .D(n2277), .Y(n1013) );
  NAND3X1 U130 ( .A(n1003), .B(n2267), .C(n2733), .Y(n1015) );
  OAI21X1 U132 ( .A(n2733), .B(n2500), .C(n1003), .Y(n1014) );
  NAND3X1 U138 ( .A(n2853), .B(n2852), .C(n2854), .Y(n1018) );
  OAI21X1 U140 ( .A(n2132), .B(n2814), .C(n2237), .Y(n1894) );
  OAI21X1 U142 ( .A(n2132), .B(n2813), .C(n2236), .Y(n1895) );
  OAI21X1 U144 ( .A(n2132), .B(n2816), .C(n2599), .Y(n1896) );
  OAI21X1 U146 ( .A(n1028), .B(n2877), .C(n2235), .Y(n1897) );
  OAI21X1 U149 ( .A(n1028), .B(n2889), .C(n2234), .Y(n1898) );
  OAI21X1 U152 ( .A(n1028), .B(n2851), .C(n2233), .Y(n1899) );
  NOR3X1 U155 ( .A(n2848), .B(reset), .C(n2775), .Y(n1028) );
  NOR3X1 U156 ( .A(n2730), .B(WE), .C(n1039), .Y(n1900) );
  NOR3X1 U157 ( .A(n2302), .B(n2421), .C(n2420), .Y(n1039) );
  NOR3X1 U160 ( .A(n1045), .B(n1046), .C(n1047), .Y(n1044) );
  XOR2X1 U161 ( .A(n2934), .B(n2613), .Y(n1047) );
  XOR2X1 U163 ( .A(n2935), .B(n2495), .Y(n1046) );
  OAI21X1 U165 ( .A(DIN[15]), .B(n2930), .C(n2142), .Y(n1045) );
  AOI22X1 U166 ( .A(n1054), .B(n2703), .C(n1055), .D(n2938), .Y(n1053) );
  OAI21X1 U167 ( .A(n2265), .B(n2275), .C(n2930), .Y(n1055) );
  NAND3X1 U168 ( .A(n2944), .B(n2943), .C(n2945), .Y(n1058) );
  NAND3X1 U169 ( .A(n2942), .B(n2941), .C(n2301), .Y(n1057) );
  NOR3X1 U172 ( .A(n2402), .B(n1066), .C(n1067), .Y(n1043) );
  XOR2X1 U173 ( .A(n2936), .B(n2524), .Y(n1067) );
  XOR2X1 U175 ( .A(n2937), .B(n2560), .Y(n1066) );
  NAND3X1 U177 ( .A(n1072), .B(n1073), .C(n1074), .Y(n1065) );
  XOR2X1 U178 ( .A(n2437), .B(n2638), .Y(n1074) );
  XOR2X1 U180 ( .A(n2485), .B(n2572), .Y(n1073) );
  XOR2X1 U182 ( .A(n2518), .B(n2708), .Y(n1072) );
  NOR3X1 U185 ( .A(n1080), .B(n1081), .C(n1082), .Y(n1079) );
  XNOR2X1 U186 ( .A(n2623), .B(n2559), .Y(n1082) );
  XNOR2X1 U188 ( .A(n2565), .B(n2461), .Y(n1081) );
  OAI21X1 U190 ( .A(DIN[15]), .B(n2880), .C(n2141), .Y(n1080) );
  AOI22X1 U191 ( .A(n1087), .B(n2716), .C(n1088), .D(n2881), .Y(n1086) );
  OAI21X1 U193 ( .A(n2395), .B(n2884), .C(n2880), .Y(n1088) );
  NOR3X1 U195 ( .A(n2581), .B(n2653), .C(n2724), .Y(n1092) );
  NAND3X1 U196 ( .A(n2883), .B(n2882), .C(n2396), .Y(n1090) );
  NOR3X1 U202 ( .A(n2401), .B(n1097), .C(n1098), .Y(n1078) );
  XNOR2X1 U203 ( .A(n2626), .B(n2670), .Y(n1098) );
  XNOR2X1 U205 ( .A(n2627), .B(n2520), .Y(n1097) );
  NAND3X1 U207 ( .A(n1101), .B(n1102), .C(n1103), .Y(n1096) );
  XOR2X1 U208 ( .A(n2422), .B(n2573), .Y(n1103) );
  XOR2X1 U210 ( .A(n2436), .B(n2529), .Y(n1102) );
  XOR2X1 U212 ( .A(n2455), .B(n2639), .Y(n1101) );
  NOR3X1 U216 ( .A(n1109), .B(n1110), .C(n1111), .Y(n1108) );
  XOR2X1 U217 ( .A(n2901), .B(n2614), .Y(n1111) );
  XOR2X1 U219 ( .A(n2900), .B(n2464), .Y(n1110) );
  OAI21X1 U221 ( .A(DIN[15]), .B(n2905), .C(n2140), .Y(n1109) );
  AOI22X1 U222 ( .A(n1118), .B(n2702), .C(n1119), .D(n2897), .Y(n1117) );
  OAI21X1 U223 ( .A(n2264), .B(n2274), .C(n2905), .Y(n1119) );
  NAND3X1 U224 ( .A(n2891), .B(n2892), .C(n2890), .Y(n1122) );
  NAND3X1 U225 ( .A(n2893), .B(n2894), .C(n2300), .Y(n1121) );
  NOR3X1 U228 ( .A(n2404), .B(n1130), .C(n1131), .Y(n1107) );
  XOR2X1 U229 ( .A(n2899), .B(n2496), .Y(n1131) );
  XOR2X1 U231 ( .A(n2898), .B(n2561), .Y(n1130) );
  NAND3X1 U233 ( .A(n1136), .B(n1137), .C(n1138), .Y(n1129) );
  XOR2X1 U234 ( .A(n2438), .B(n2636), .Y(n1138) );
  XOR2X1 U236 ( .A(n2457), .B(n2706), .Y(n1137) );
  XOR2X1 U238 ( .A(n2487), .B(n2570), .Y(n1136) );
  NOR3X1 U241 ( .A(n1144), .B(n1145), .C(n1146), .Y(n1143) );
  XNOR2X1 U242 ( .A(n2624), .B(n2492), .Y(n1146) );
  XNOR2X1 U244 ( .A(n2566), .B(n2462), .Y(n1145) );
  OAI21X1 U246 ( .A(DIN[15]), .B(n2949), .C(n2139), .Y(n1144) );
  AOI22X1 U247 ( .A(n1151), .B(n2717), .C(n1152), .D(n2950), .Y(n1150) );
  OAI21X1 U249 ( .A(n2397), .B(n2953), .C(n2949), .Y(n1152) );
  NOR3X1 U251 ( .A(n2582), .B(n2654), .C(n2725), .Y(n1156) );
  NAND3X1 U252 ( .A(n2952), .B(n2951), .C(n2398), .Y(n1154) );
  NOR3X1 U258 ( .A(n2403), .B(n1161), .C(n1162), .Y(n1142) );
  XNOR2X1 U259 ( .A(n2628), .B(n2671), .Y(n1162) );
  XNOR2X1 U261 ( .A(n2629), .B(n2521), .Y(n1161) );
  NAND3X1 U263 ( .A(n1165), .B(n1166), .C(n1167), .Y(n1160) );
  XOR2X1 U264 ( .A(n2423), .B(n2574), .Y(n1167) );
  XOR2X1 U266 ( .A(n2456), .B(n2530), .Y(n1166) );
  XOR2X1 U268 ( .A(n2486), .B(n2640), .Y(n1165) );
  NAND3X1 U270 ( .A(n2468), .B(n2527), .C(n2299), .Y(n1040) );
  NOR3X1 U273 ( .A(n1174), .B(n1175), .C(n1176), .Y(n1173) );
  XOR2X1 U274 ( .A(n2858), .B(n2497), .Y(n1176) );
  XOR2X1 U276 ( .A(n2862), .B(n2562), .Y(n1175) );
  OAI21X1 U278 ( .A(DIN[11]), .B(n2859), .C(n2138), .Y(n1174) );
  AOI22X1 U279 ( .A(n1183), .B(n2701), .C(n1184), .D(n2867), .Y(n1182) );
  OAI21X1 U280 ( .A(n2263), .B(n2273), .C(n2859), .Y(n1184) );
  NAND3X1 U281 ( .A(n2869), .B(n2868), .C(n2870), .Y(n1187) );
  NAND3X1 U282 ( .A(n2866), .B(n2865), .C(n2298), .Y(n1186) );
  NOR3X1 U285 ( .A(n2435), .B(n1195), .C(n1196), .Y(n1172) );
  XOR2X1 U286 ( .A(n2861), .B(n2616), .Y(n1196) );
  XOR2X1 U288 ( .A(n2860), .B(n2465), .Y(n1195) );
  NAND3X1 U290 ( .A(n1201), .B(n1202), .C(n1203), .Y(n1194) );
  XOR2X1 U291 ( .A(n2458), .B(n2569), .Y(n1203) );
  XOR2X1 U293 ( .A(n2519), .B(n2705), .Y(n1202) );
  XOR2X1 U295 ( .A(n2488), .B(n2635), .Y(n1201) );
  NOR3X1 U298 ( .A(n1209), .B(n1210), .C(n1211), .Y(n1208) );
  XNOR2X1 U299 ( .A(n2632), .B(n2672), .Y(n1211) );
  XNOR2X1 U301 ( .A(n2633), .B(n2493), .Y(n1210) );
  OAI21X1 U303 ( .A(DIN[11]), .B(n2963), .C(n2137), .Y(n1209) );
  AOI22X1 U304 ( .A(n1216), .B(n2718), .C(n1217), .D(n2966), .Y(n1215) );
  OAI21X1 U306 ( .A(n2416), .B(n2967), .C(n2963), .Y(n1217) );
  NOR3X1 U308 ( .A(n2584), .B(n2656), .C(n2727), .Y(n1221) );
  NAND3X1 U309 ( .A(n2965), .B(n2964), .C(n2417), .Y(n1219) );
  NOR3X1 U315 ( .A(n2419), .B(n1226), .C(n1227), .Y(n1207) );
  XNOR2X1 U316 ( .A(n2634), .B(n2523), .Y(n1227) );
  XNOR2X1 U318 ( .A(n2568), .B(n2463), .Y(n1226) );
  NAND3X1 U320 ( .A(n1230), .B(n1231), .C(n1232), .Y(n1225) );
  XOR2X1 U321 ( .A(n2439), .B(n2532), .Y(n1232) );
  XOR2X1 U323 ( .A(n2459), .B(n2642), .Y(n1231) );
  XOR2X1 U325 ( .A(n2489), .B(n2576), .Y(n1230) );
  NOR3X1 U328 ( .A(n1238), .B(n1239), .C(n1240), .Y(n1237) );
  XOR2X1 U329 ( .A(n2920), .B(n2615), .Y(n1240) );
  XOR2X1 U331 ( .A(n2919), .B(n2466), .Y(n1239) );
  OAI21X1 U333 ( .A(DIN[15]), .B(n2924), .C(n2136), .Y(n1238) );
  AOI22X1 U334 ( .A(n1247), .B(n2704), .C(n1248), .D(n2916), .Y(n1246) );
  OAI21X1 U335 ( .A(n2262), .B(n2272), .C(n2924), .Y(n1248) );
  NAND3X1 U336 ( .A(n2910), .B(n2911), .C(n2909), .Y(n1251) );
  NAND3X1 U337 ( .A(n2912), .B(n2913), .C(n2297), .Y(n1250) );
  NOR3X1 U340 ( .A(n2418), .B(n1259), .C(n1260), .Y(n1236) );
  XOR2X1 U341 ( .A(n2918), .B(n2498), .Y(n1260) );
  XOR2X1 U343 ( .A(n2917), .B(n2563), .Y(n1259) );
  NAND3X1 U345 ( .A(n1265), .B(n1266), .C(n1267), .Y(n1258) );
  XOR2X1 U346 ( .A(n2441), .B(n2637), .Y(n1267) );
  XOR2X1 U348 ( .A(n2460), .B(n2707), .Y(n1266) );
  XOR2X1 U350 ( .A(n2491), .B(n2571), .Y(n1265) );
  NOR3X1 U353 ( .A(n1273), .B(n1274), .C(n1275), .Y(n1272) );
  XNOR2X1 U354 ( .A(n2625), .B(n2494), .Y(n1275) );
  XNOR2X1 U356 ( .A(n2567), .B(n2442), .Y(n1274) );
  OAI21X1 U358 ( .A(DIN[15]), .B(n2956), .C(n2135), .Y(n1273) );
  AOI22X1 U359 ( .A(n1280), .B(n2719), .C(n1281), .D(n2957), .Y(n1279) );
  OAI21X1 U361 ( .A(n2399), .B(n2960), .C(n2956), .Y(n1281) );
  NOR3X1 U363 ( .A(n2583), .B(n2655), .C(n2726), .Y(n1285) );
  NAND3X1 U364 ( .A(n2959), .B(n2958), .C(n2400), .Y(n1283) );
  NOR3X1 U370 ( .A(n2405), .B(n1290), .C(n1291), .Y(n1271) );
  XNOR2X1 U371 ( .A(n2630), .B(n2673), .Y(n1291) );
  XNOR2X1 U373 ( .A(n2631), .B(n2522), .Y(n1290) );
  NAND3X1 U375 ( .A(n1294), .B(n1295), .C(n1296), .Y(n1289) );
  XOR2X1 U376 ( .A(n2424), .B(n2575), .Y(n1296) );
  XOR2X1 U378 ( .A(n2440), .B(n2531), .Y(n1295) );
  XOR2X1 U380 ( .A(n2490), .B(n2641), .Y(n1294) );
  OAI21X1 U382 ( .A(n2132), .B(n2743), .C(n2232), .Y(n1901) );
  OAI21X1 U384 ( .A(n2132), .B(n2745), .C(n2231), .Y(n1902) );
  OAI21X1 U386 ( .A(n2132), .B(n2746), .C(n2445), .Y(n1903) );
  OAI21X1 U388 ( .A(n2132), .B(n2744), .C(n2230), .Y(n1904) );
  OAI21X1 U390 ( .A(n2132), .B(n2739), .C(n2229), .Y(n1905) );
  OAI21X1 U392 ( .A(n2132), .B(n2740), .C(n2387), .Y(n1906) );
  OAI21X1 U394 ( .A(n2132), .B(n2741), .C(n2228), .Y(n1907) );
  OAI21X1 U396 ( .A(n2132), .B(n2742), .C(n2227), .Y(n1908) );
  OAI21X1 U398 ( .A(n2132), .B(n2817), .C(n2473), .Y(n1909) );
  OAI21X1 U400 ( .A(n2132), .B(n2819), .C(n2545), .Y(n1910) );
  OAI21X1 U402 ( .A(n2132), .B(n2820), .C(n2505), .Y(n1911) );
  OAI21X1 U404 ( .A(n2132), .B(n2821), .C(n2226), .Y(n1912) );
  OAI21X1 U406 ( .A(n2132), .B(n2822), .C(n2225), .Y(n1913) );
  OAI21X1 U408 ( .A(n2132), .B(n2824), .C(n2407), .Y(n1914) );
  OAI21X1 U410 ( .A(n2132), .B(n2825), .C(n2427), .Y(n1915) );
  OAI21X1 U412 ( .A(n2132), .B(n2826), .C(n2446), .Y(n1916) );
  NAND3X1 U414 ( .A(n2846), .B(n2847), .C(n2544), .Y(n1021) );
  OAI21X1 U415 ( .A(n1335), .B(n2928), .C(n2224), .Y(n1917) );
  OAI21X1 U418 ( .A(n1335), .B(n2929), .C(n2223), .Y(n1918) );
  OAI21X1 U421 ( .A(n1335), .B(n2309), .C(n2669), .Y(n1919) );
  OAI21X1 U424 ( .A(n1335), .B(n2930), .C(n2222), .Y(n1920) );
  OAI21X1 U427 ( .A(n1335), .B(n2931), .C(n2517), .Y(n1921) );
  OAI21X1 U430 ( .A(n1335), .B(n2932), .C(n2554), .Y(n1922) );
  OAI21X1 U433 ( .A(n1335), .B(n2933), .C(n2608), .Y(n1923) );
  OAI21X1 U436 ( .A(n1335), .B(n2934), .C(n2221), .Y(n1924) );
  OAI21X1 U439 ( .A(n1335), .B(n2935), .C(n2220), .Y(n1925) );
  OAI21X1 U442 ( .A(n1335), .B(n2936), .C(n2219), .Y(n1926) );
  OAI21X1 U445 ( .A(n1335), .B(n2937), .C(n2218), .Y(n1927) );
  OAI21X1 U448 ( .A(n1335), .B(n2938), .C(n2391), .Y(n1928) );
  OAI21X1 U451 ( .A(n1335), .B(n2939), .C(n2555), .Y(n1929) );
  OAI21X1 U454 ( .A(n1335), .B(n2940), .C(n2609), .Y(n1930) );
  OAI21X1 U457 ( .A(n1335), .B(n2941), .C(n2410), .Y(n1931) );
  OAI21X1 U460 ( .A(n1335), .B(n2942), .C(n2430), .Y(n1932) );
  OAI21X1 U463 ( .A(n1335), .B(n2943), .C(n2450), .Y(n1933) );
  OAI21X1 U466 ( .A(n1335), .B(n2944), .C(n2476), .Y(n1934) );
  OAI21X1 U469 ( .A(n1335), .B(n2945), .C(n2506), .Y(n1935) );
  NOR3X1 U472 ( .A(n2747), .B(n2665), .C(n2594), .Y(n1335) );
  OAI21X1 U473 ( .A(n2814), .B(n2131), .C(n2217), .Y(n1936) );
  OAI21X1 U475 ( .A(n2813), .B(n2131), .C(n2216), .Y(n1937) );
  OAI21X1 U477 ( .A(n2816), .B(n2131), .C(n2215), .Y(n1938) );
  OAI21X1 U479 ( .A(n2743), .B(n2131), .C(n2214), .Y(n1939) );
  OAI21X1 U481 ( .A(n2745), .B(n2131), .C(n2213), .Y(n1940) );
  OAI21X1 U483 ( .A(n2746), .B(n2131), .C(n2507), .Y(n1941) );
  OAI21X1 U485 ( .A(n2744), .B(n2131), .C(n2212), .Y(n1942) );
  OAI21X1 U487 ( .A(n2739), .B(n2131), .C(n2211), .Y(n1943) );
  OAI21X1 U489 ( .A(n2740), .B(n2131), .C(n2411), .Y(n1944) );
  OAI21X1 U491 ( .A(n2741), .B(n2131), .C(n2392), .Y(n1945) );
  OAI21X1 U493 ( .A(n2742), .B(n2131), .C(n2210), .Y(n1946) );
  OAI21X1 U495 ( .A(n2817), .B(n2131), .C(n2600), .Y(n1947) );
  OAI21X1 U497 ( .A(n2819), .B(n2131), .C(n2431), .Y(n1948) );
  OAI21X1 U499 ( .A(n2820), .B(n2131), .C(n2546), .Y(n1949) );
  OAI21X1 U501 ( .A(n2821), .B(n2131), .C(n2209), .Y(n1950) );
  OAI21X1 U503 ( .A(n2822), .B(n2131), .C(n2208), .Y(n1951) );
  OAI21X1 U505 ( .A(n2824), .B(n2131), .C(n2508), .Y(n1952) );
  OAI21X1 U507 ( .A(n2825), .B(n2131), .C(n2451), .Y(n1953) );
  OAI21X1 U509 ( .A(n2826), .B(n2131), .C(n2477), .Y(n1954) );
  NAND3X1 U511 ( .A(n2544), .B(n2846), .C(n2665), .Y(n1371) );
  OAI21X1 U512 ( .A(n1391), .B(n2908), .C(n2428), .Y(n1955) );
  OAI21X1 U515 ( .A(n1391), .B(n2907), .C(n2408), .Y(n1956) );
  OAI21X1 U518 ( .A(n1391), .B(n2906), .C(n2514), .Y(n1957) );
  OAI21X1 U521 ( .A(n1391), .B(n2905), .C(n2389), .Y(n1958) );
  OAI21X1 U524 ( .A(n1391), .B(n2904), .C(n2552), .Y(n1959) );
  OAI21X1 U527 ( .A(n1391), .B(n2903), .C(n2483), .Y(n1960) );
  OAI21X1 U530 ( .A(n1391), .B(n2902), .C(n2454), .Y(n1961) );
  OAI21X1 U533 ( .A(n1391), .B(n2901), .C(n2448), .Y(n1962) );
  OAI21X1 U536 ( .A(n1391), .B(n2900), .C(n2207), .Y(n1963) );
  OAI21X1 U539 ( .A(n1391), .B(n2899), .C(n2206), .Y(n1964) );
  OAI21X1 U542 ( .A(n1391), .B(n2898), .C(n2205), .Y(n1965) );
  OAI21X1 U545 ( .A(n1391), .B(n2897), .C(n2204), .Y(n1966) );
  OAI21X1 U548 ( .A(n1391), .B(n2896), .C(n2551), .Y(n1967) );
  OAI21X1 U551 ( .A(n1391), .B(n2895), .C(n2605), .Y(n1968) );
  OAI21X1 U554 ( .A(n1391), .B(n2894), .C(n2474), .Y(n1969) );
  OAI21X1 U557 ( .A(n1391), .B(n2893), .C(n2203), .Y(n1970) );
  OAI21X1 U560 ( .A(n1391), .B(n2892), .C(n2202), .Y(n1971) );
  OAI21X1 U563 ( .A(n1391), .B(n2891), .C(n2201), .Y(n1972) );
  OAI21X1 U566 ( .A(n1391), .B(n2890), .C(n2200), .Y(n1973) );
  NOR3X1 U569 ( .A(n2594), .B(n2747), .C(n2847), .Y(n1391) );
  OAI21X1 U570 ( .A(n2814), .B(n2130), .C(n2199), .Y(n1974) );
  OAI21X1 U572 ( .A(n2813), .B(n2130), .C(n2198), .Y(n1975) );
  OAI21X1 U574 ( .A(n2816), .B(n2130), .C(n2197), .Y(n1976) );
  OAI21X1 U576 ( .A(n2743), .B(n2130), .C(n2196), .Y(n1977) );
  OAI21X1 U578 ( .A(n2745), .B(n2130), .C(n2195), .Y(n1978) );
  OAI21X1 U580 ( .A(n2746), .B(n2130), .C(n2478), .Y(n1979) );
  OAI21X1 U582 ( .A(n2744), .B(n2130), .C(n2194), .Y(n1980) );
  OAI21X1 U584 ( .A(n2739), .B(n2130), .C(n2193), .Y(n1981) );
  OAI21X1 U586 ( .A(n2740), .B(n2130), .C(n2192), .Y(n1982) );
  OAI21X1 U588 ( .A(n2741), .B(n2130), .C(n2412), .Y(n1983) );
  OAI21X1 U590 ( .A(n2742), .B(n2130), .C(n2393), .Y(n1984) );
  OAI21X1 U592 ( .A(n2817), .B(n2130), .C(n2432), .Y(n1985) );
  OAI21X1 U594 ( .A(n2819), .B(n2130), .C(n2452), .Y(n1986) );
  OAI21X1 U596 ( .A(n2820), .B(n2130), .C(n2601), .Y(n1987) );
  OAI21X1 U598 ( .A(n2821), .B(n2130), .C(n2191), .Y(n1988) );
  OAI21X1 U600 ( .A(n2822), .B(n2130), .C(n2190), .Y(n1989) );
  OAI21X1 U602 ( .A(n2824), .B(n2130), .C(n2479), .Y(n1990) );
  OAI21X1 U604 ( .A(n2825), .B(n2130), .C(n2509), .Y(n1991) );
  OAI21X1 U606 ( .A(n2826), .B(n2130), .C(n2547), .Y(n1992) );
  NAND3X1 U608 ( .A(n2544), .B(n2847), .C(n2747), .Y(n1417) );
  OAI21X1 U609 ( .A(n1437), .B(n2927), .C(n2449), .Y(n1993) );
  OAI21X1 U612 ( .A(n1437), .B(n2926), .C(n2668), .Y(n1994) );
  OAI21X1 U615 ( .A(n1437), .B(n2925), .C(n2553), .Y(n1995) );
  OAI21X1 U618 ( .A(n1437), .B(n2924), .C(n2429), .Y(n1996) );
  OAI21X1 U621 ( .A(n1437), .B(n2923), .C(n2607), .Y(n1997) );
  OAI21X1 U624 ( .A(n1437), .B(n2922), .C(n2516), .Y(n1998) );
  OAI21X1 U627 ( .A(n1437), .B(n2921), .C(n2484), .Y(n1999) );
  OAI21X1 U630 ( .A(n1437), .B(n2920), .C(n2475), .Y(n2000) );
  OAI21X1 U633 ( .A(n1437), .B(n2919), .C(n2409), .Y(n2001) );
  OAI21X1 U636 ( .A(n1437), .B(n2918), .C(n2390), .Y(n2002) );
  OAI21X1 U639 ( .A(n1437), .B(n2917), .C(n2189), .Y(n2003) );
  OAI21X1 U642 ( .A(n1437), .B(n2916), .C(n2188), .Y(n2004) );
  OAI21X1 U645 ( .A(n1437), .B(n2915), .C(n2515), .Y(n2005) );
  OAI21X1 U648 ( .A(n1437), .B(n2914), .C(n2606), .Y(n2006) );
  OAI21X1 U651 ( .A(n1437), .B(n2913), .C(n2187), .Y(n2007) );
  OAI21X1 U654 ( .A(n1437), .B(n2912), .C(n2186), .Y(n2008) );
  OAI21X1 U657 ( .A(n1437), .B(n2911), .C(n2185), .Y(n2009) );
  OAI21X1 U660 ( .A(n1437), .B(n2910), .C(n2184), .Y(n2010) );
  OAI21X1 U663 ( .A(n1437), .B(n2909), .C(n2183), .Y(n2011) );
  NOR3X1 U666 ( .A(n2594), .B(n2665), .C(n2846), .Y(n1437) );
  OAI21X1 U667 ( .A(n2814), .B(n2129), .C(n2182), .Y(n2012) );
  OAI21X1 U670 ( .A(n2813), .B(n2129), .C(n2181), .Y(n2013) );
  OAI21X1 U673 ( .A(n2816), .B(n2129), .C(n2180), .Y(n2014) );
  OAI21X1 U676 ( .A(n2743), .B(n2129), .C(n2179), .Y(n2015) );
  OAI21X1 U678 ( .A(n2745), .B(n2129), .C(n2510), .Y(n2016) );
  OAI21X1 U680 ( .A(n2746), .B(n2129), .C(n2548), .Y(n2017) );
  OAI21X1 U682 ( .A(n2744), .B(n2129), .C(n2178), .Y(n2018) );
  OAI21X1 U684 ( .A(n2739), .B(n2129), .C(n2177), .Y(n2019) );
  OAI21X1 U686 ( .A(n2740), .B(n2129), .C(n2176), .Y(n2020) );
  OAI21X1 U688 ( .A(n2741), .B(n2129), .C(n2175), .Y(n2021) );
  OAI21X1 U690 ( .A(n2742), .B(n2129), .C(n2413), .Y(n2022) );
  OAI21X1 U692 ( .A(n2817), .B(n2129), .C(n2174), .Y(n2023) );
  OAI21X1 U695 ( .A(n2819), .B(n2129), .C(n2394), .Y(n2024) );
  OAI21X1 U698 ( .A(n2820), .B(n2129), .C(n2433), .Y(n2025) );
  OAI21X1 U701 ( .A(n2821), .B(n2129), .C(n2453), .Y(n2026) );
  OAI21X1 U704 ( .A(n2822), .B(n2129), .C(n2511), .Y(n2027) );
  OAI21X1 U707 ( .A(n2824), .B(n2129), .C(n2549), .Y(n2028) );
  OAI21X1 U710 ( .A(n2825), .B(n2129), .C(n2480), .Y(n2029) );
  OAI21X1 U713 ( .A(n2826), .B(n2129), .C(n2602), .Y(n2030) );
  NAND3X1 U715 ( .A(n2665), .B(n2544), .C(n2747), .Y(n1463) );
  AOI21X1 U716 ( .A(n2469), .B(n2873), .C(n2776), .Y(n1334) );
  OAI21X1 U718 ( .A(n1485), .B(n2852), .C(n2173), .Y(n2031) );
  OAI21X1 U721 ( .A(n1485), .B(n2853), .C(n2172), .Y(n2032) );
  OAI21X1 U724 ( .A(n1485), .B(n2854), .C(n2171), .Y(n2033) );
  OAI21X1 U727 ( .A(n1485), .B(n2855), .C(n2513), .Y(n2034) );
  OAI21X1 U732 ( .A(n1485), .B(n2856), .C(n2482), .Y(n2035) );
  OAI21X1 U737 ( .A(n1485), .B(n2857), .C(n2603), .Y(n2036) );
  OAI21X1 U742 ( .A(n1485), .B(n2858), .C(n2425), .Y(n2037) );
  OAI21X1 U747 ( .A(n1485), .B(n2859), .C(n2170), .Y(n2038) );
  OAI21X1 U752 ( .A(n1485), .B(n2860), .C(n2169), .Y(n2039) );
  OAI21X1 U757 ( .A(n1485), .B(n2861), .C(n2168), .Y(n2040) );
  OAI21X1 U762 ( .A(n1485), .B(n2862), .C(n2167), .Y(n2041) );
  OAI21X1 U767 ( .A(n1485), .B(n2863), .C(n2550), .Y(n2042) );
  OAI21X1 U770 ( .A(n1485), .B(n2864), .C(n2604), .Y(n2043) );
  OAI21X1 U773 ( .A(n1485), .B(n2865), .C(n2166), .Y(n2044) );
  OAI21X1 U776 ( .A(n1485), .B(n2866), .C(n2386), .Y(n2045) );
  OAI21X1 U779 ( .A(n1485), .B(n2867), .C(n2406), .Y(n2046) );
  OAI21X1 U782 ( .A(n1485), .B(n2868), .C(n2426), .Y(n2047) );
  OAI21X1 U785 ( .A(n1485), .B(n2869), .C(n2444), .Y(n2048) );
  OAI21X1 U788 ( .A(n1485), .B(n2870), .C(n2472), .Y(n2049) );
  NOR3X1 U791 ( .A(n2847), .B(n2594), .C(n2846), .Y(n1485) );
  AOI21X1 U793 ( .A(n2848), .B(last[2]), .C(n2382), .Y(n1368) );
  OAI21X1 U798 ( .A(n2874), .B(n2271), .C(n2540), .Y(n1037) );
  AOI21X1 U799 ( .A(n1514), .B(n2385), .C(n2383), .Y(n1512) );
  OAI21X1 U801 ( .A(n2304), .B(n2353), .C(n2307), .Y(n1514) );
  AOI21X1 U805 ( .A(n2848), .B(last[1]), .C(n2308), .Y(n1369) );
  NAND3X1 U806 ( .A(n2503), .B(n2540), .C(n2286), .Y(n1034) );
  NAND3X1 U807 ( .A(n2385), .B(n2384), .C(n2351), .Y(n1523) );
  NAND3X1 U809 ( .A(n2248), .B(n2353), .C(n2296), .Y(n1525) );
  NAND3X1 U812 ( .A(n2661), .B(n2738), .C(n2590), .Y(n1520) );
  NAND3X1 U813 ( .A(n2593), .B(n2737), .C(n2657), .Y(n1521) );
  NAND3X1 U814 ( .A(n2385), .B(n2384), .C(n1528), .Y(n1031) );
  NAND3X1 U816 ( .A(n2658), .B(n2734), .C(n2587), .Y(n1513) );
  NAND3X1 U817 ( .A(n2731), .B(n2663), .C(n2541), .Y(n1522) );
  NAND3X1 U818 ( .A(n2732), .B(n2664), .C(n2542), .Y(n1517) );
  NAND3X1 U819 ( .A(n2659), .B(n2735), .C(n2588), .Y(n1515) );
  NAND3X1 U820 ( .A(n2660), .B(n2736), .C(n2589), .Y(n1519) );
  NAND3X1 U821 ( .A(n2543), .B(n2596), .C(n2504), .Y(n1526) );
  OAI21X1 U822 ( .A(n2831), .B(n2969), .C(n2159), .Y(n2050) );
  NAND3X1 U823 ( .A(n2734), .B(n2969), .C(n2830), .Y(n1531) );
  OAI21X1 U825 ( .A(n2734), .B(n1534), .C(n1535), .Y(n2051) );
  OAI21X1 U827 ( .A(n2261), .B(n2872), .C(n2158), .Y(n2052) );
  NAND3X1 U828 ( .A(n2842), .B(n2731), .C(n2295), .Y(n1540) );
  AOI21X1 U830 ( .A(n2842), .B(n2876), .C(n1545), .Y(n1538) );
  OAI21X1 U831 ( .A(n2843), .B(n2876), .C(n2157), .Y(n2053) );
  NAND3X1 U832 ( .A(n2663), .B(n2876), .C(n2842), .Y(n1547) );
  OAI21X1 U835 ( .A(n2663), .B(n1548), .C(n2379), .Y(n1545) );
  OAI21X1 U836 ( .A(n2663), .B(n1548), .C(n1550), .Y(n2054) );
  OAI21X1 U838 ( .A(n2946), .B(n2340), .C(n2379), .Y(n1548) );
  NAND3X1 U841 ( .A(n85), .B(n2871), .C(n1556), .Y(n1553) );
  NAND3X1 U845 ( .A(n2350), .B(n2875), .C(n2285), .Y(n1558) );
  AOI21X1 U846 ( .A(n2731), .B(n2773), .C(n89), .Y(n1561) );
  NAND3X1 U848 ( .A(n2350), .B(n2876), .C(n88), .Y(n1557) );
  OAI21X1 U851 ( .A(n2260), .B(n2886), .C(n2156), .Y(n2055) );
  NAND3X1 U852 ( .A(n2840), .B(n2732), .C(n2294), .Y(n1567) );
  AOI21X1 U854 ( .A(n2840), .B(n2888), .C(n1572), .Y(n1565) );
  OAI21X1 U855 ( .A(n2841), .B(n2888), .C(n2155), .Y(n2056) );
  NAND3X1 U856 ( .A(n2664), .B(n2888), .C(n2840), .Y(n1574) );
  OAI21X1 U859 ( .A(n2664), .B(n1575), .C(n2376), .Y(n1572) );
  OAI21X1 U860 ( .A(n2664), .B(n1575), .C(n1577), .Y(n2057) );
  OAI21X1 U862 ( .A(n2946), .B(n2336), .C(n2376), .Y(n1575) );
  NAND3X1 U865 ( .A(n84), .B(n2968), .C(n1556), .Y(n1579) );
  NAND3X1 U869 ( .A(n2349), .B(n2887), .C(n2284), .Y(n1582) );
  AOI21X1 U870 ( .A(n2732), .B(n2773), .C(n89), .Y(n1585) );
  NAND3X1 U872 ( .A(n2349), .B(n2888), .C(n88), .Y(n1581) );
  OAI21X1 U875 ( .A(n2259), .B(n2972), .C(n2154), .Y(n2058) );
  NAND3X1 U876 ( .A(n2838), .B(n2659), .C(n2293), .Y(n1588) );
  AOI21X1 U878 ( .A(n2838), .B(n2974), .C(n1593), .Y(n1586) );
  OAI21X1 U879 ( .A(n2839), .B(n2974), .C(n2153), .Y(n2059) );
  NAND3X1 U880 ( .A(n2735), .B(n2974), .C(n2838), .Y(n1595) );
  OAI21X1 U883 ( .A(n2735), .B(n1596), .C(n2372), .Y(n1593) );
  OAI21X1 U884 ( .A(n2735), .B(n1596), .C(n1598), .Y(n2060) );
  OAI21X1 U886 ( .A(n2946), .B(n2332), .C(n2372), .Y(n1596) );
  NAND3X1 U889 ( .A(n2871), .B(n2968), .C(n1556), .Y(n1600) );
  NAND3X1 U893 ( .A(n2348), .B(n2973), .C(n2283), .Y(n1603) );
  AOI21X1 U894 ( .A(n2659), .B(n2773), .C(n89), .Y(n1606) );
  NAND3X1 U896 ( .A(n2348), .B(n2974), .C(n88), .Y(n1602) );
  OAI21X1 U899 ( .A(n2258), .B(n2978), .C(n2152), .Y(n2061) );
  NAND3X1 U900 ( .A(n2836), .B(n2661), .C(n2292), .Y(n1609) );
  AOI21X1 U902 ( .A(n2836), .B(n2980), .C(n1614), .Y(n1607) );
  OAI21X1 U903 ( .A(n2837), .B(n2980), .C(n2151), .Y(n2062) );
  NAND3X1 U904 ( .A(n2738), .B(n2980), .C(n2836), .Y(n1616) );
  OAI21X1 U907 ( .A(n2738), .B(n1617), .C(n2369), .Y(n1614) );
  OAI21X1 U908 ( .A(n2738), .B(n1617), .C(n1619), .Y(n2063) );
  OAI21X1 U910 ( .A(n2946), .B(n2328), .C(n2369), .Y(n1617) );
  NAND3X1 U913 ( .A(n85), .B(n84), .C(n1623), .Y(n1621) );
  NAND3X1 U917 ( .A(n2347), .B(n2979), .C(n2282), .Y(n1625) );
  AOI21X1 U918 ( .A(n2661), .B(n2773), .C(n89), .Y(n1628) );
  NAND3X1 U920 ( .A(n2347), .B(n2980), .C(n88), .Y(n1624) );
  OAI21X1 U923 ( .A(n2257), .B(n2975), .C(n2150), .Y(n2064) );
  NAND3X1 U924 ( .A(n2834), .B(n2593), .C(n2291), .Y(n1631) );
  AOI21X1 U926 ( .A(n2834), .B(n2977), .C(n1636), .Y(n1629) );
  OAI21X1 U927 ( .A(n2835), .B(n2977), .C(n2149), .Y(n2065) );
  NAND3X1 U928 ( .A(n2737), .B(n2977), .C(n2834), .Y(n1638) );
  OAI21X1 U931 ( .A(n2737), .B(n1639), .C(n2366), .Y(n1636) );
  OAI21X1 U932 ( .A(n2737), .B(n1639), .C(n1641), .Y(n2066) );
  OAI21X1 U934 ( .A(n2946), .B(n2324), .C(n2366), .Y(n1639) );
  NAND3X1 U937 ( .A(n85), .B(n2871), .C(n1623), .Y(n1643) );
  NAND3X1 U941 ( .A(n2564), .B(n2976), .C(n2281), .Y(n1646) );
  AOI21X1 U942 ( .A(n2593), .B(n2773), .C(n89), .Y(n1649) );
  NAND3X1 U944 ( .A(n2564), .B(n2977), .C(n88), .Y(n1645) );
  OAI21X1 U947 ( .A(n2256), .B(n2981), .C(n2148), .Y(n2067) );
  NAND3X1 U948 ( .A(n2832), .B(n2660), .C(n2290), .Y(n1652) );
  AOI21X1 U950 ( .A(n2832), .B(n2983), .C(n1657), .Y(n1650) );
  OAI21X1 U951 ( .A(n2833), .B(n2983), .C(n2147), .Y(n2068) );
  NAND3X1 U952 ( .A(n2736), .B(n2983), .C(n2832), .Y(n1659) );
  OAI21X1 U955 ( .A(n2736), .B(n1660), .C(n2362), .Y(n1657) );
  OAI21X1 U956 ( .A(n2736), .B(n1660), .C(n1662), .Y(n2069) );
  OAI21X1 U958 ( .A(n2946), .B(n2320), .C(n2362), .Y(n1660) );
  NAND3X1 U961 ( .A(n84), .B(n2968), .C(n1623), .Y(n1664) );
  NAND3X1 U965 ( .A(n2346), .B(n2982), .C(n2280), .Y(n1667) );
  AOI21X1 U966 ( .A(n2660), .B(n2773), .C(n89), .Y(n1670) );
  NAND3X1 U968 ( .A(n2346), .B(n2983), .C(n88), .Y(n1666) );
  OAI21X1 U971 ( .A(n2255), .B(n2850), .C(n2146), .Y(n2070) );
  NAND3X1 U972 ( .A(n2828), .B(n2543), .C(n2289), .Y(n1673) );
  AOI21X1 U974 ( .A(n2828), .B(n2849), .C(n1678), .Y(n1671) );
  OAI21X1 U975 ( .A(n2829), .B(n2849), .C(n2145), .Y(n2071) );
  NAND3X1 U976 ( .A(n2596), .B(n2849), .C(n2828), .Y(n1680) );
  OAI21X1 U979 ( .A(n2596), .B(n1681), .C(n2354), .Y(n1678) );
  OAI21X1 U980 ( .A(n2254), .B(n2971), .C(n2144), .Y(n2072) );
  NAND3X1 U981 ( .A(n2830), .B(n2658), .C(n2288), .Y(n1685) );
  AOI21X1 U983 ( .A(n2830), .B(n2969), .C(n1533), .Y(n1683) );
  OAI21X1 U984 ( .A(n2734), .B(n1534), .C(n2358), .Y(n1533) );
  OAI21X1 U986 ( .A(n2946), .B(n2316), .C(n2358), .Y(n1534) );
  NAND3X1 U989 ( .A(n85), .B(n84), .C(n1556), .Y(n1688) );
  NOR3X1 U990 ( .A(n2752), .B(j_3_), .C(n2885), .Y(n1556) );
  NAND3X1 U995 ( .A(n2345), .B(n2970), .C(n2279), .Y(n1691) );
  AOI21X1 U996 ( .A(n2658), .B(n2773), .C(n89), .Y(n1694) );
  NAND3X1 U998 ( .A(n2345), .B(n2969), .C(n88), .Y(n1690) );
  OAI21X1 U1001 ( .A(n2596), .B(n1681), .C(n1695), .Y(n2073) );
  OAI21X1 U1003 ( .A(n2946), .B(n2312), .C(n2354), .Y(n1681) );
  NAND3X1 U1010 ( .A(n2871), .B(n2968), .C(n1623), .Y(n1697) );
  NOR3X1 U1011 ( .A(j_3_), .B(n86), .C(n2752), .Y(n1623) );
  NAND3X1 U1018 ( .A(n2344), .B(n2845), .C(n2278), .Y(n1700) );
  AOI21X1 U1019 ( .A(n2543), .B(n2773), .C(n89), .Y(n1703) );
  NAND3X1 U1023 ( .A(n2344), .B(n2849), .C(n88), .Y(n1699) );
  AND2X1 U1209 ( .A(n2534), .B(DIN[12]), .Y(n1212) );
  AND2X1 U1210 ( .A(n2582), .B(DIN[9]), .Y(n1163) );
  AND2X1 U1211 ( .A(n2581), .B(DIN[9]), .Y(n1099) );
  AND2X1 U1212 ( .A(n2533), .B(DIN[11]), .Y(n1083) );
  AND2X1 U1213 ( .A(n2583), .B(DIN[9]), .Y(n1292) );
  AND2X1 U1214 ( .A(n2305), .B(n2307), .Y(n1524) );
  AND2X1 U1215 ( .A(n2591), .B(n2537), .Y(n905) );
  OR2X1 U1216 ( .A(n2362), .B(n2982), .Y(n1662) );
  OR2X1 U1217 ( .A(n2369), .B(n2979), .Y(n1619) );
  OR2X1 U1218 ( .A(n2366), .B(n2976), .Y(n1641) );
  OR2X1 U1219 ( .A(n2372), .B(n2973), .Y(n1598) );
  OR2X1 U1220 ( .A(n2358), .B(n2970), .Y(n1535) );
  AND2X1 U1221 ( .A(n2752), .B(n2557), .Y(n1781) );
  AND2X1 U1222 ( .A(match), .B(n2827), .Y(n874) );
  OR2X1 U1223 ( .A(n2376), .B(n2887), .Y(n1577) );
  OR2X1 U1224 ( .A(n2379), .B(n2875), .Y(n1550) );
  OR2X1 U1225 ( .A(n2354), .B(n2845), .Y(n1695) );
  OR2X1 U1226 ( .A(n2844), .B(n2730), .Y(n904) );
  AND2X1 U1227 ( .A(n2617), .B(EN), .Y(n868) );
  AND2X1 U1228 ( .A(n1017), .B(n2538), .Y(n1003) );
  AND2X1 U1229 ( .A(n2503), .B(n2540), .Y(n1528) );
  OR2X1 U1230 ( .A(n2666), .B(WE), .Y(n878) );
  BUFX2 U1231 ( .A(n921), .Y(n2074) );
  BUFX2 U1232 ( .A(mem[104]), .Y(n2075) );
  BUFX2 U1233 ( .A(mem[105]), .Y(n2076) );
  BUFX2 U1234 ( .A(mem[106]), .Y(n2077) );
  BUFX2 U1235 ( .A(mem[107]), .Y(n2078) );
  BUFX2 U1236 ( .A(mem[111]), .Y(n2079) );
  BUFX2 U1237 ( .A(matchN[19]), .Y(n2080) );
  BUFX2 U1238 ( .A(matchN[20]), .Y(n2081) );
  BUFX2 U1239 ( .A(matchN[8]), .Y(n2082) );
  BUFX2 U1240 ( .A(matchN[7]), .Y(n2083) );
  BUFX2 U1241 ( .A(mem[47]), .Y(n2084) );
  BUFX2 U1242 ( .A(mem[43]), .Y(n2085) );
  BUFX2 U1243 ( .A(mem[42]), .Y(n2086) );
  BUFX2 U1244 ( .A(mem[41]), .Y(n2087) );
  BUFX2 U1245 ( .A(mem[40]), .Y(n2088) );
  BUFX2 U1246 ( .A(matchN[14]), .Y(n2089) );
  BUFX2 U1247 ( .A(matchN[13]), .Y(n2090) );
  BUFX2 U1248 ( .A(mem[79]), .Y(n2091) );
  BUFX2 U1249 ( .A(mem[75]), .Y(n2092) );
  BUFX2 U1250 ( .A(mem[74]), .Y(n2093) );
  BUFX2 U1251 ( .A(mem[73]), .Y(n2094) );
  BUFX2 U1252 ( .A(mem[72]), .Y(n2095) );
  BUFX2 U1253 ( .A(mem[8]), .Y(n2096) );
  BUFX2 U1254 ( .A(mem[9]), .Y(n2097) );
  BUFX2 U1255 ( .A(mem[10]), .Y(n2098) );
  BUFX2 U1256 ( .A(mem[11]), .Y(n2099) );
  BUFX2 U1257 ( .A(mem[12]), .Y(n2100) );
  BUFX2 U1258 ( .A(n2990), .Y(n2101) );
  BUFX2 U1259 ( .A(n2993), .Y(n2102) );
  BUFX2 U1260 ( .A(n2996), .Y(n2103) );
  BUFX2 U1261 ( .A(n1699), .Y(n2104) );
  BUFX2 U1262 ( .A(n1700), .Y(n2105) );
  BUFX2 U1263 ( .A(n1697), .Y(n2106) );
  BUFX2 U1264 ( .A(n1690), .Y(n2107) );
  BUFX2 U1265 ( .A(n1691), .Y(n2108) );
  BUFX2 U1266 ( .A(n1688), .Y(n2109) );
  BUFX2 U1267 ( .A(n1666), .Y(n2110) );
  BUFX2 U1268 ( .A(n1667), .Y(n2111) );
  BUFX2 U1269 ( .A(n1664), .Y(n2112) );
  BUFX2 U1270 ( .A(n1645), .Y(n2113) );
  BUFX2 U1271 ( .A(n1646), .Y(n2114) );
  BUFX2 U1272 ( .A(n1643), .Y(n2115) );
  BUFX2 U1273 ( .A(n1624), .Y(n2116) );
  BUFX2 U1274 ( .A(n1625), .Y(n2117) );
  BUFX2 U1275 ( .A(n1621), .Y(n2118) );
  BUFX2 U1276 ( .A(n1602), .Y(n2119) );
  BUFX2 U1277 ( .A(n1603), .Y(n2120) );
  BUFX2 U1278 ( .A(n1600), .Y(n2121) );
  BUFX2 U1279 ( .A(n1581), .Y(n2122) );
  BUFX2 U1280 ( .A(n1582), .Y(n2123) );
  BUFX2 U1281 ( .A(n1579), .Y(n2124) );
  BUFX2 U1282 ( .A(n1557), .Y(n2125) );
  BUFX2 U1283 ( .A(n1558), .Y(n2126) );
  BUFX2 U1284 ( .A(n1553), .Y(n2127) );
  BUFX2 U1285 ( .A(n1525), .Y(n2128) );
  BUFX2 U1286 ( .A(n1463), .Y(n2129) );
  BUFX2 U1287 ( .A(n1417), .Y(n2130) );
  BUFX2 U1288 ( .A(n1371), .Y(n2131) );
  BUFX2 U1289 ( .A(n1021), .Y(n2132) );
  BUFX2 U1290 ( .A(n908), .Y(n2133) );
  BUFX2 U1291 ( .A(n882), .Y(n2134) );
  OR2X1 U1292 ( .A(n2314), .B(n2315), .Y(n2312) );
  OR2X1 U1293 ( .A(n1701), .B(n2313), .Y(n2315) );
  OR2X1 U1294 ( .A(n2318), .B(n2319), .Y(n2316) );
  OR2X1 U1295 ( .A(n1692), .B(n2317), .Y(n2319) );
  OR2X1 U1296 ( .A(n2322), .B(n2323), .Y(n2320) );
  OR2X1 U1297 ( .A(n1668), .B(n2321), .Y(n2323) );
  OR2X1 U1298 ( .A(n2326), .B(n2327), .Y(n2324) );
  OR2X1 U1299 ( .A(n1647), .B(n2325), .Y(n2327) );
  OR2X1 U1300 ( .A(n2330), .B(n2331), .Y(n2328) );
  OR2X1 U1301 ( .A(n1626), .B(n2329), .Y(n2331) );
  OR2X1 U1302 ( .A(n2334), .B(n2335), .Y(n2332) );
  OR2X1 U1303 ( .A(n1604), .B(n2333), .Y(n2335) );
  OR2X1 U1304 ( .A(n2338), .B(n2339), .Y(n2336) );
  OR2X1 U1305 ( .A(n1583), .B(n2337), .Y(n2339) );
  OR2X1 U1306 ( .A(n2342), .B(n2343), .Y(n2340) );
  OR2X1 U1307 ( .A(n1559), .B(n2341), .Y(n2343) );
  OR2X1 U1308 ( .A(n2356), .B(n2357), .Y(n2354) );
  OR2X1 U1309 ( .A(n1698), .B(n2355), .Y(n2357) );
  OR2X1 U1310 ( .A(n2360), .B(n2361), .Y(n2358) );
  OR2X1 U1311 ( .A(n1689), .B(n2359), .Y(n2361) );
  OR2X1 U1312 ( .A(n2364), .B(n2365), .Y(n2362) );
  OR2X1 U1313 ( .A(n1665), .B(n2363), .Y(n2365) );
  OR2X1 U1314 ( .A(n2367), .B(n2368), .Y(n2366) );
  OR2X1 U1315 ( .A(n1644), .B(n2359), .Y(n2368) );
  OR2X1 U1316 ( .A(n2370), .B(n2371), .Y(n2369) );
  OR2X1 U1317 ( .A(n1622), .B(n2355), .Y(n2371) );
  OR2X1 U1318 ( .A(n2374), .B(n2375), .Y(n2372) );
  OR2X1 U1319 ( .A(n1601), .B(n2373), .Y(n2375) );
  OR2X1 U1320 ( .A(n2377), .B(n2378), .Y(n2376) );
  OR2X1 U1321 ( .A(n1580), .B(n2363), .Y(n2378) );
  OR2X1 U1322 ( .A(n2380), .B(n2381), .Y(n2379) );
  OR2X1 U1323 ( .A(n1554), .B(n2373), .Y(n2381) );
  AND2X1 U1324 ( .A(n2818), .B(n2815), .Y(n2989) );
  AND2X1 U1325 ( .A(n87), .B(n2850), .Y(n1701) );
  AND2X1 U1326 ( .A(n868), .B(n2312), .Y(n1698) );
  AND2X1 U1327 ( .A(n87), .B(n2971), .Y(n1692) );
  AND2X1 U1328 ( .A(n868), .B(n2316), .Y(n1689) );
  AND2X1 U1329 ( .A(n87), .B(n2981), .Y(n1668) );
  AND2X1 U1330 ( .A(n868), .B(n2320), .Y(n1665) );
  AND2X1 U1331 ( .A(n87), .B(n2975), .Y(n1647) );
  AND2X1 U1332 ( .A(n868), .B(n2324), .Y(n1644) );
  AND2X1 U1333 ( .A(n87), .B(n2978), .Y(n1626) );
  AND2X1 U1334 ( .A(n868), .B(n2328), .Y(n1622) );
  AND2X1 U1335 ( .A(n87), .B(n2972), .Y(n1604) );
  AND2X1 U1336 ( .A(n868), .B(n2332), .Y(n1601) );
  AND2X1 U1337 ( .A(n87), .B(n2886), .Y(n1583) );
  AND2X1 U1338 ( .A(n868), .B(n2336), .Y(n1580) );
  AND2X1 U1339 ( .A(n87), .B(n2872), .Y(n1559) );
  AND2X1 U1340 ( .A(n868), .B(n2340), .Y(n1554) );
  BUFX2 U1341 ( .A(n1279), .Y(n2135) );
  BUFX2 U1342 ( .A(n1246), .Y(n2136) );
  BUFX2 U1343 ( .A(n1215), .Y(n2137) );
  BUFX2 U1344 ( .A(n1182), .Y(n2138) );
  BUFX2 U1345 ( .A(n1150), .Y(n2139) );
  BUFX2 U1346 ( .A(n1117), .Y(n2140) );
  BUFX2 U1347 ( .A(n1086), .Y(n2141) );
  BUFX2 U1348 ( .A(n1053), .Y(n2142) );
  BUFX2 U1349 ( .A(n1013), .Y(n2143) );
  BUFX2 U1350 ( .A(n1685), .Y(n2144) );
  BUFX2 U1351 ( .A(n1680), .Y(n2145) );
  BUFX2 U1352 ( .A(n1673), .Y(n2146) );
  BUFX2 U1353 ( .A(n1659), .Y(n2147) );
  BUFX2 U1354 ( .A(n1652), .Y(n2148) );
  BUFX2 U1355 ( .A(n1638), .Y(n2149) );
  BUFX2 U1356 ( .A(n1631), .Y(n2150) );
  BUFX2 U1357 ( .A(n1616), .Y(n2151) );
  BUFX2 U1358 ( .A(n1609), .Y(n2152) );
  BUFX2 U1359 ( .A(n1595), .Y(n2153) );
  BUFX2 U1360 ( .A(n1588), .Y(n2154) );
  BUFX2 U1361 ( .A(n1574), .Y(n2155) );
  BUFX2 U1362 ( .A(n1567), .Y(n2156) );
  BUFX2 U1363 ( .A(n1547), .Y(n2157) );
  BUFX2 U1364 ( .A(n1540), .Y(n2158) );
  BUFX2 U1365 ( .A(n1531), .Y(n2159) );
  BUFX2 U1366 ( .A(n1007), .Y(n2160) );
  BUFX2 U1367 ( .A(n1000), .Y(n2161) );
  BUFX2 U1368 ( .A(n985), .Y(n2162) );
  BUFX2 U1369 ( .A(n969), .Y(n2163) );
  BUFX2 U1370 ( .A(n954), .Y(n2164) );
  BUFX2 U1371 ( .A(n938), .Y(n2165) );
  AND2X1 U1372 ( .A(n1485), .B(DIN[5]), .Y(n1504) );
  INVX1 U1373 ( .A(n1504), .Y(n2166) );
  AND2X1 U1374 ( .A(n1485), .B(n1314), .Y(n1499) );
  INVX1 U1375 ( .A(n1499), .Y(n2167) );
  AND2X1 U1376 ( .A(n1485), .B(n1312), .Y(n1498) );
  INVX1 U1377 ( .A(n1498), .Y(n2168) );
  AND2X1 U1378 ( .A(n1485), .B(n1310), .Y(n1497) );
  INVX1 U1379 ( .A(n1497), .Y(n2169) );
  AND2X1 U1380 ( .A(n1485), .B(n1308), .Y(n1496) );
  INVX1 U1381 ( .A(n1496), .Y(n2170) );
  AND2X1 U1382 ( .A(n1485), .B(n250), .Y(n1488) );
  INVX1 U1383 ( .A(n1488), .Y(n2171) );
  AND2X1 U1384 ( .A(n1485), .B(n251), .Y(n1487) );
  INVX1 U1385 ( .A(n1487), .Y(n2172) );
  AND2X1 U1386 ( .A(n1485), .B(n252), .Y(n1486) );
  INVX1 U1387 ( .A(n1486), .Y(n2173) );
  AND2X1 U1388 ( .A(n2650), .B(n2129), .Y(n1475) );
  INVX1 U1389 ( .A(n1475), .Y(n2174) );
  AND2X1 U1390 ( .A(n2634), .B(n2129), .Y(n1473) );
  INVX1 U1391 ( .A(n1473), .Y(n2175) );
  AND2X1 U1392 ( .A(n2568), .B(n2129), .Y(n1472) );
  INVX1 U1393 ( .A(n1472), .Y(n2176) );
  AND2X1 U1394 ( .A(n2620), .B(n2129), .Y(n1471) );
  INVX1 U1395 ( .A(n1471), .Y(n2177) );
  AND2X1 U1396 ( .A(n2632), .B(n2129), .Y(n1470) );
  INVX1 U1397 ( .A(n1470), .Y(n2178) );
  AND2X1 U1398 ( .A(n2532), .B(n2129), .Y(n1467) );
  INVX1 U1399 ( .A(n1467), .Y(n2179) );
  AND2X1 U1400 ( .A(n2662), .B(n2129), .Y(n1466) );
  INVX1 U1401 ( .A(n1466), .Y(n2180) );
  AND2X1 U1402 ( .A(n2539), .B(n2129), .Y(n1465) );
  INVX1 U1403 ( .A(n1465), .Y(n2181) );
  AND2X1 U1404 ( .A(n2715), .B(n2129), .Y(n1464) );
  INVX1 U1405 ( .A(n1464), .Y(n2182) );
  AND2X1 U1406 ( .A(n1437), .B(DIN[0]), .Y(n1462) );
  INVX1 U1407 ( .A(n1462), .Y(n2183) );
  AND2X1 U1408 ( .A(n1437), .B(DIN[1]), .Y(n1461) );
  INVX1 U1409 ( .A(n1461), .Y(n2184) );
  AND2X1 U1410 ( .A(n1437), .B(DIN[2]), .Y(n1460) );
  INVX1 U1411 ( .A(n1460), .Y(n2185) );
  AND2X1 U1412 ( .A(n1437), .B(DIN[3]), .Y(n1459) );
  INVX1 U1413 ( .A(n1459), .Y(n2186) );
  AND2X1 U1414 ( .A(n1437), .B(DIN[4]), .Y(n1458) );
  INVX1 U1415 ( .A(n1458), .Y(n2187) );
  AND2X1 U1416 ( .A(n1437), .B(DIN[7]), .Y(n1453) );
  INVX1 U1417 ( .A(n1453), .Y(n2188) );
  AND2X1 U1418 ( .A(n1437), .B(n1314), .Y(n1452) );
  INVX1 U1419 ( .A(n1452), .Y(n2189) );
  AND2X1 U1420 ( .A(n2536), .B(n2130), .Y(n1433) );
  INVX1 U1421 ( .A(n1433), .Y(n2190) );
  AND2X1 U1422 ( .A(n2579), .B(n2130), .Y(n1432) );
  INVX1 U1423 ( .A(n1432), .Y(n2191) );
  AND2X1 U1424 ( .A(n2567), .B(n2130), .Y(n1426) );
  INVX1 U1425 ( .A(n1426), .Y(n2192) );
  AND2X1 U1426 ( .A(n2625), .B(n2130), .Y(n1425) );
  INVX1 U1427 ( .A(n1425), .Y(n2193) );
  AND2X1 U1428 ( .A(n2641), .B(n2130), .Y(n1424) );
  INVX1 U1429 ( .A(n1424), .Y(n2194) );
  AND2X1 U1430 ( .A(n2531), .B(n2130), .Y(n1422) );
  INVX1 U1431 ( .A(n1422), .Y(n2195) );
  AND2X1 U1432 ( .A(n2621), .B(n2130), .Y(n1421) );
  INVX1 U1433 ( .A(n1421), .Y(n2196) );
  AND2X1 U1434 ( .A(n2729), .B(n2130), .Y(n1420) );
  INVX1 U1435 ( .A(n1420), .Y(n2197) );
  AND2X1 U1436 ( .A(n2691), .B(n2130), .Y(n1419) );
  INVX1 U1437 ( .A(n1419), .Y(n2198) );
  AND2X1 U1438 ( .A(n2714), .B(n2130), .Y(n1418) );
  INVX1 U1439 ( .A(n1418), .Y(n2199) );
  AND2X1 U1440 ( .A(n1391), .B(DIN[0]), .Y(n1416) );
  INVX1 U1441 ( .A(n1416), .Y(n2200) );
  AND2X1 U1442 ( .A(n1391), .B(DIN[1]), .Y(n1415) );
  INVX1 U1443 ( .A(n1415), .Y(n2201) );
  AND2X1 U1444 ( .A(n1391), .B(DIN[2]), .Y(n1414) );
  INVX1 U1445 ( .A(n1414), .Y(n2202) );
  AND2X1 U1446 ( .A(n1391), .B(DIN[3]), .Y(n1413) );
  INVX1 U1447 ( .A(n1413), .Y(n2203) );
  AND2X1 U1448 ( .A(n1391), .B(DIN[7]), .Y(n1407) );
  INVX1 U1449 ( .A(n1407), .Y(n2204) );
  AND2X1 U1450 ( .A(n1391), .B(n1314), .Y(n1406) );
  INVX1 U1451 ( .A(n1406), .Y(n2205) );
  AND2X1 U1452 ( .A(n1391), .B(n1312), .Y(n1405) );
  INVX1 U1453 ( .A(n1405), .Y(n2206) );
  AND2X1 U1454 ( .A(n1391), .B(n1310), .Y(n1404) );
  INVX1 U1455 ( .A(n1404), .Y(n2207) );
  AND2X1 U1456 ( .A(n2535), .B(n2131), .Y(n1387) );
  INVX1 U1457 ( .A(n1387), .Y(n2208) );
  AND2X1 U1458 ( .A(n2578), .B(n2131), .Y(n1386) );
  INVX1 U1459 ( .A(n1386), .Y(n2209) );
  AND2X1 U1460 ( .A(n2629), .B(n2131), .Y(n1382) );
  INVX1 U1461 ( .A(n1382), .Y(n2210) );
  AND2X1 U1462 ( .A(n2624), .B(n2131), .Y(n1379) );
  INVX1 U1463 ( .A(n1379), .Y(n2211) );
  AND2X1 U1464 ( .A(n2640), .B(n2131), .Y(n1378) );
  INVX1 U1465 ( .A(n1378), .Y(n2212) );
  AND2X1 U1466 ( .A(n2530), .B(n2131), .Y(n1376) );
  INVX1 U1467 ( .A(n1376), .Y(n2213) );
  AND2X1 U1468 ( .A(n2619), .B(n2131), .Y(n1375) );
  INVX1 U1469 ( .A(n1375), .Y(n2214) );
  AND2X1 U1470 ( .A(n2728), .B(n2131), .Y(n1374) );
  INVX1 U1471 ( .A(n1374), .Y(n2215) );
  AND2X1 U1472 ( .A(n2690), .B(n2131), .Y(n1373) );
  INVX1 U1473 ( .A(n1373), .Y(n2216) );
  AND2X1 U1474 ( .A(n2713), .B(n2131), .Y(n1372) );
  INVX1 U1475 ( .A(n1372), .Y(n2217) );
  AND2X1 U1476 ( .A(n1335), .B(n1314), .Y(n1356) );
  INVX1 U1477 ( .A(n1356), .Y(n2218) );
  AND2X1 U1478 ( .A(n1335), .B(n1312), .Y(n1354) );
  INVX1 U1479 ( .A(n1354), .Y(n2219) );
  AND2X1 U1480 ( .A(n1335), .B(n1310), .Y(n1352) );
  INVX1 U1481 ( .A(n1352), .Y(n2220) );
  AND2X1 U1482 ( .A(n1335), .B(n1308), .Y(n1350) );
  INVX1 U1483 ( .A(n1350), .Y(n2221) );
  AND2X1 U1484 ( .A(n1335), .B(n1300), .Y(n1339) );
  INVX1 U1485 ( .A(n1339), .Y(n2222) );
  AND2X1 U1486 ( .A(n1335), .B(n251), .Y(n1337) );
  INVX1 U1487 ( .A(n1337), .Y(n2223) );
  AND2X1 U1488 ( .A(n1335), .B(n252), .Y(n1336) );
  INVX1 U1489 ( .A(n1336), .Y(n2224) );
  AND2X1 U1490 ( .A(n2533), .B(n2132), .Y(n1325) );
  INVX1 U1491 ( .A(n1325), .Y(n2225) );
  AND2X1 U1492 ( .A(n2577), .B(n2132), .Y(n1323) );
  INVX1 U1493 ( .A(n1323), .Y(n2226) );
  AND2X1 U1494 ( .A(n2627), .B(n2132), .Y(n1315) );
  INVX1 U1495 ( .A(n1315), .Y(n2227) );
  AND2X1 U1496 ( .A(n2626), .B(n2132), .Y(n1313) );
  INVX1 U1497 ( .A(n1313), .Y(n2228) );
  AND2X1 U1498 ( .A(n2623), .B(n2132), .Y(n1309) );
  INVX1 U1499 ( .A(n1309), .Y(n2229) );
  AND2X1 U1500 ( .A(n2639), .B(n2132), .Y(n1307) );
  INVX1 U1501 ( .A(n1307), .Y(n2230) );
  AND2X1 U1502 ( .A(n2529), .B(n2132), .Y(n1303) );
  INVX1 U1503 ( .A(n1303), .Y(n2231) );
  AND2X1 U1504 ( .A(n2618), .B(n2132), .Y(n1301) );
  INVX1 U1505 ( .A(n1301), .Y(n2232) );
  AND2X1 U1506 ( .A(n1028), .B(n1037), .Y(n1036) );
  INVX1 U1507 ( .A(n1036), .Y(n2233) );
  AND2X1 U1508 ( .A(n1028), .B(n2308), .Y(n1033) );
  INVX1 U1509 ( .A(n1033), .Y(n2234) );
  AND2X1 U1510 ( .A(n1028), .B(n2382), .Y(n1030) );
  INVX1 U1511 ( .A(n1030), .Y(n2235) );
  AND2X1 U1512 ( .A(n2694), .B(n2132), .Y(n1025) );
  INVX1 U1513 ( .A(n1025), .Y(n2236) );
  AND2X1 U1514 ( .A(n2693), .B(n2132), .Y(n1023) );
  INVX1 U1515 ( .A(n1023), .Y(n2237) );
  AND2X1 U1516 ( .A(n2750), .B(n991), .Y(n990) );
  INVX1 U1517 ( .A(n990), .Y(n2238) );
  AND2X1 U1518 ( .A(n2471), .B(n2750), .Y(n987) );
  INVX1 U1519 ( .A(n987), .Y(n2239) );
  AND2X1 U1520 ( .A(n2585), .B(n975), .Y(n974) );
  INVX1 U1521 ( .A(n974), .Y(n2240) );
  AND2X1 U1522 ( .A(n2753), .B(n960), .Y(n959) );
  INVX1 U1523 ( .A(n959), .Y(n2241) );
  AND2X1 U1524 ( .A(n2311), .B(n2753), .Y(n956) );
  INVX1 U1525 ( .A(n956), .Y(n2242) );
  AND2X1 U1526 ( .A(n2597), .B(n944), .Y(n943) );
  INVX1 U1527 ( .A(n943), .Y(n2243) );
  AND2X1 U1528 ( .A(n2748), .B(n926), .Y(n925) );
  INVX1 U1529 ( .A(n925), .Y(n2244) );
  BUFX2 U1530 ( .A(n883), .Y(n2245) );
  OR2X1 U1531 ( .A(n972), .B(n2808), .Y(n971) );
  INVX1 U1532 ( .A(n971), .Y(n2246) );
  OR2X1 U1533 ( .A(n941), .B(n2804), .Y(n940) );
  INVX1 U1534 ( .A(n940), .Y(n2247) );
  BUFX2 U1535 ( .A(n1526), .Y(n2248) );
  BUFX2 U1536 ( .A(n909), .Y(n2249) );
  AND2X1 U1537 ( .A(n2955), .B(n975), .Y(n986) );
  INVX1 U1538 ( .A(n986), .Y(n2250) );
  AND2X1 U1539 ( .A(n2948), .B(n944), .Y(n955) );
  INVX1 U1540 ( .A(n955), .Y(n2251) );
  AND2X1 U1541 ( .A(n2799), .B(n2700), .Y(n915) );
  INVX1 U1542 ( .A(n915), .Y(n2252) );
  BUFX2 U1543 ( .A(n884), .Y(n2253) );
  BUFX2 U1544 ( .A(n1683), .Y(n2254) );
  BUFX2 U1545 ( .A(n1671), .Y(n2255) );
  BUFX2 U1546 ( .A(n1650), .Y(n2256) );
  BUFX2 U1547 ( .A(n1629), .Y(n2257) );
  BUFX2 U1548 ( .A(n1607), .Y(n2258) );
  BUFX2 U1549 ( .A(n1586), .Y(n2259) );
  BUFX2 U1550 ( .A(n1565), .Y(n2260) );
  BUFX2 U1551 ( .A(n1538), .Y(n2261) );
  BUFX2 U1552 ( .A(n1250), .Y(n2262) );
  BUFX2 U1553 ( .A(n1186), .Y(n2263) );
  BUFX2 U1554 ( .A(n1121), .Y(n2264) );
  BUFX2 U1555 ( .A(n1057), .Y(n2265) );
  BUFX2 U1556 ( .A(n910), .Y(n2266) );
  AND2X1 U1557 ( .A(n2662), .B(n2854), .Y(n1016) );
  INVX1 U1558 ( .A(n1016), .Y(n2267) );
  AND2X1 U1559 ( .A(n2926), .B(n991), .Y(n1001) );
  INVX1 U1560 ( .A(n1001), .Y(n2268) );
  AND2X1 U1561 ( .A(n2907), .B(n960), .Y(n970) );
  INVX1 U1562 ( .A(n970), .Y(n2269) );
  AND2X1 U1563 ( .A(n2929), .B(n926), .Y(n939) );
  INVX1 U1564 ( .A(n939), .Y(n2270) );
  BUFX2 U1565 ( .A(n1512), .Y(n2271) );
  BUFX2 U1566 ( .A(n1251), .Y(n2272) );
  BUFX2 U1567 ( .A(n1187), .Y(n2273) );
  BUFX2 U1568 ( .A(n1122), .Y(n2274) );
  BUFX2 U1569 ( .A(n1058), .Y(n2275) );
  BUFX2 U1570 ( .A(n895), .Y(n2276) );
  BUFX2 U1571 ( .A(n1015), .Y(n2277) );
  BUFX2 U1572 ( .A(n1703), .Y(n2278) );
  BUFX2 U1573 ( .A(n1694), .Y(n2279) );
  BUFX2 U1574 ( .A(n1670), .Y(n2280) );
  BUFX2 U1575 ( .A(n1649), .Y(n2281) );
  BUFX2 U1576 ( .A(n1628), .Y(n2282) );
  BUFX2 U1577 ( .A(n1606), .Y(n2283) );
  BUFX2 U1578 ( .A(n1585), .Y(n2284) );
  BUFX2 U1579 ( .A(n1561), .Y(n2285) );
  BUFX2 U1580 ( .A(n1523), .Y(n2286) );
  BUFX2 U1581 ( .A(n911), .Y(n2287) );
  OR2X1 U1582 ( .A(n2587), .B(n2970), .Y(n1686) );
  INVX1 U1583 ( .A(n1686), .Y(n2288) );
  OR2X1 U1584 ( .A(n2504), .B(n2845), .Y(n1675) );
  INVX1 U1585 ( .A(n1675), .Y(n2289) );
  OR2X1 U1586 ( .A(n2589), .B(n2982), .Y(n1654) );
  INVX1 U1587 ( .A(n1654), .Y(n2290) );
  OR2X1 U1588 ( .A(n2657), .B(n2976), .Y(n1633) );
  INVX1 U1589 ( .A(n1633), .Y(n2291) );
  OR2X1 U1590 ( .A(n2590), .B(n2979), .Y(n1611) );
  INVX1 U1591 ( .A(n1611), .Y(n2292) );
  OR2X1 U1592 ( .A(n2588), .B(n2973), .Y(n1590) );
  INVX1 U1593 ( .A(n1590), .Y(n2293) );
  OR2X1 U1594 ( .A(n2542), .B(n2887), .Y(n1569) );
  INVX1 U1595 ( .A(n1569), .Y(n2294) );
  OR2X1 U1596 ( .A(n2541), .B(n2875), .Y(n1542) );
  INVX1 U1597 ( .A(n1542), .Y(n2295) );
  OR2X1 U1598 ( .A(n2382), .B(n2351), .Y(n1527) );
  INVX1 U1599 ( .A(n1527), .Y(n2296) );
  OR2X1 U1600 ( .A(n2646), .B(n2712), .Y(n1257) );
  INVX1 U1601 ( .A(n1257), .Y(n2297) );
  OR2X1 U1602 ( .A(n2643), .B(n2709), .Y(n1193) );
  INVX1 U1603 ( .A(n1193), .Y(n2298) );
  OR2X1 U1604 ( .A(n1011), .B(n1017), .Y(n1171) );
  INVX1 U1605 ( .A(n1171), .Y(n2299) );
  OR2X1 U1606 ( .A(n2644), .B(n2710), .Y(n1128) );
  INVX1 U1607 ( .A(n1128), .Y(n2300) );
  OR2X1 U1608 ( .A(n2645), .B(n2711), .Y(n1064) );
  INVX1 U1609 ( .A(n1064), .Y(n2301) );
  BUFX2 U1610 ( .A(n1040), .Y(n2302) );
  BUFX2 U1611 ( .A(n2999), .Y(match) );
  INVX1 U1612 ( .A(n2305), .Y(n2304) );
  BUFX2 U1613 ( .A(n1521), .Y(n2305) );
  BUFX2 U1614 ( .A(n928), .Y(n2306) );
  BUFX2 U1615 ( .A(n1520), .Y(n2307) );
  BUFX2 U1616 ( .A(n1034), .Y(n2308) );
  INVX1 U1617 ( .A(n2310), .Y(n2309) );
  BUFX2 U1618 ( .A(matchN[18]), .Y(n2310) );
  BUFX2 U1619 ( .A(n957), .Y(n2311) );
  INVX1 U1620 ( .A(n2105), .Y(n2313) );
  INVX1 U1621 ( .A(n2104), .Y(n2314) );
  INVX1 U1622 ( .A(n2108), .Y(n2317) );
  INVX1 U1623 ( .A(n2107), .Y(n2318) );
  INVX1 U1624 ( .A(n2111), .Y(n2321) );
  INVX1 U1625 ( .A(n2110), .Y(n2322) );
  INVX1 U1626 ( .A(n2114), .Y(n2325) );
  INVX1 U1627 ( .A(n2113), .Y(n2326) );
  INVX1 U1628 ( .A(n2117), .Y(n2329) );
  INVX1 U1629 ( .A(n2116), .Y(n2330) );
  INVX1 U1630 ( .A(n2120), .Y(n2333) );
  INVX1 U1631 ( .A(n2119), .Y(n2334) );
  INVX1 U1632 ( .A(n2123), .Y(n2337) );
  INVX1 U1633 ( .A(n2122), .Y(n2338) );
  INVX1 U1634 ( .A(n2126), .Y(n2341) );
  INVX1 U1635 ( .A(n2125), .Y(n2342) );
  AND2X1 U1636 ( .A(n2504), .B(n2774), .Y(n1702) );
  INVX1 U1637 ( .A(n1702), .Y(n2344) );
  AND2X1 U1638 ( .A(n2587), .B(n2774), .Y(n1693) );
  INVX1 U1639 ( .A(n1693), .Y(n2345) );
  AND2X1 U1640 ( .A(n2589), .B(n2774), .Y(n1669) );
  INVX1 U1641 ( .A(n1669), .Y(n2346) );
  AND2X1 U1642 ( .A(n2590), .B(n2774), .Y(n1627) );
  INVX1 U1643 ( .A(n1627), .Y(n2347) );
  AND2X1 U1644 ( .A(n2588), .B(n2774), .Y(n1605) );
  INVX1 U1645 ( .A(n1605), .Y(n2348) );
  AND2X1 U1646 ( .A(n2542), .B(n2774), .Y(n1584) );
  INVX1 U1647 ( .A(n1584), .Y(n2349) );
  AND2X1 U1648 ( .A(n2541), .B(n2774), .Y(n1560) );
  INVX1 U1649 ( .A(n1560), .Y(n2350) );
  INVX1 U1650 ( .A(n1524), .Y(n2351) );
  BUFX2 U1651 ( .A(n923), .Y(n2352) );
  BUFX2 U1652 ( .A(n1519), .Y(n2353) );
  INVX1 U1653 ( .A(n2775), .Y(n2355) );
  INVX1 U1654 ( .A(n2106), .Y(n2356) );
  INVX1 U1655 ( .A(n2775), .Y(n2359) );
  INVX1 U1656 ( .A(n2109), .Y(n2360) );
  INVX1 U1657 ( .A(n2775), .Y(n2363) );
  INVX1 U1658 ( .A(n2112), .Y(n2364) );
  INVX1 U1659 ( .A(n2115), .Y(n2367) );
  INVX1 U1660 ( .A(n2118), .Y(n2370) );
  INVX1 U1661 ( .A(n2776), .Y(n2373) );
  INVX1 U1662 ( .A(n2121), .Y(n2374) );
  INVX1 U1663 ( .A(n2124), .Y(n2377) );
  INVX1 U1664 ( .A(n2127), .Y(n2380) );
  BUFX2 U1665 ( .A(n1031), .Y(n2382) );
  INVX1 U1666 ( .A(n2384), .Y(n2383) );
  BUFX2 U1667 ( .A(n1517), .Y(n2384) );
  BUFX2 U1668 ( .A(n1515), .Y(n2385) );
  AND2X1 U1669 ( .A(n1485), .B(DIN[4]), .Y(n1505) );
  INVX1 U1670 ( .A(n1505), .Y(n2386) );
  AND2X1 U1671 ( .A(n2565), .B(n2132), .Y(n1311) );
  INVX1 U1672 ( .A(n1311), .Y(n2387) );
  AND2X1 U1673 ( .A(n86), .B(n2666), .Y(n879) );
  INVX1 U1674 ( .A(n879), .Y(n2388) );
  AND2X1 U1675 ( .A(n1391), .B(n1300), .Y(n1396) );
  INVX1 U1676 ( .A(n1396), .Y(n2389) );
  AND2X1 U1677 ( .A(n1437), .B(n1312), .Y(n1451) );
  INVX1 U1678 ( .A(n1451), .Y(n2390) );
  AND2X1 U1679 ( .A(n1335), .B(DIN[7]), .Y(n1358) );
  INVX1 U1680 ( .A(n1358), .Y(n2391) );
  AND2X1 U1681 ( .A(n2628), .B(n2131), .Y(n1381) );
  INVX1 U1682 ( .A(n1381), .Y(n2392) );
  AND2X1 U1683 ( .A(n2631), .B(n2130), .Y(n1428) );
  INVX1 U1684 ( .A(n1428), .Y(n2393) );
  AND2X1 U1685 ( .A(n2723), .B(n2129), .Y(n1476) );
  INVX1 U1686 ( .A(n1476), .Y(n2394) );
  BUFX2 U1687 ( .A(n1090), .Y(n2395) );
  OR2X1 U1688 ( .A(n2647), .B(n2720), .Y(n1095) );
  INVX1 U1689 ( .A(n1095), .Y(n2396) );
  BUFX2 U1690 ( .A(n1154), .Y(n2397) );
  OR2X1 U1691 ( .A(n2648), .B(n2721), .Y(n1159) );
  INVX1 U1692 ( .A(n1159), .Y(n2398) );
  BUFX2 U1693 ( .A(n1283), .Y(n2399) );
  OR2X1 U1694 ( .A(n2649), .B(n2722), .Y(n1288) );
  INVX1 U1695 ( .A(n1288), .Y(n2400) );
  BUFX2 U1696 ( .A(n1096), .Y(n2401) );
  BUFX2 U1697 ( .A(n1065), .Y(n2402) );
  BUFX2 U1698 ( .A(n1160), .Y(n2403) );
  BUFX2 U1699 ( .A(n1129), .Y(n2404) );
  BUFX2 U1700 ( .A(n1289), .Y(n2405) );
  AND2X1 U1701 ( .A(n1485), .B(DIN[3]), .Y(n1506) );
  INVX1 U1702 ( .A(n1506), .Y(n2406) );
  AND2X1 U1703 ( .A(n2653), .B(n2132), .Y(n1327) );
  INVX1 U1704 ( .A(n1327), .Y(n2407) );
  AND2X1 U1705 ( .A(n1391), .B(n251), .Y(n1393) );
  INVX1 U1706 ( .A(n1393), .Y(n2408) );
  AND2X1 U1707 ( .A(n1437), .B(n1310), .Y(n1450) );
  INVX1 U1708 ( .A(n1450), .Y(n2409) );
  AND2X1 U1709 ( .A(n1335), .B(DIN[4]), .Y(n1363) );
  INVX1 U1710 ( .A(n1363), .Y(n2410) );
  AND2X1 U1711 ( .A(n2566), .B(n2131), .Y(n1380) );
  INVX1 U1712 ( .A(n1380), .Y(n2411) );
  AND2X1 U1713 ( .A(n2630), .B(n2130), .Y(n1427) );
  INVX1 U1714 ( .A(n1427), .Y(n2412) );
  AND2X1 U1715 ( .A(n2633), .B(n2129), .Y(n1474) );
  INVX1 U1716 ( .A(n1474), .Y(n2413) );
  BUFX2 U1717 ( .A(n889), .Y(n2414) );
  AND2X1 U1718 ( .A(n84), .B(n2666), .Y(n890) );
  INVX1 U1719 ( .A(n890), .Y(n2415) );
  BUFX2 U1720 ( .A(n1219), .Y(n2416) );
  OR2X1 U1721 ( .A(n2650), .B(n2723), .Y(n1224) );
  INVX1 U1722 ( .A(n1224), .Y(n2417) );
  BUFX2 U1723 ( .A(n1258), .Y(n2418) );
  BUFX2 U1724 ( .A(n1225), .Y(n2419) );
  AND2X1 U1725 ( .A(n2501), .B(n2467), .Y(n1042) );
  INVX1 U1726 ( .A(n1042), .Y(n2420) );
  AND2X1 U1727 ( .A(n2443), .B(n2526), .Y(n1041) );
  INVX1 U1728 ( .A(n1041), .Y(n2421) );
  AND2X1 U1729 ( .A(n2720), .B(DIN[13]), .Y(n1104) );
  INVX1 U1730 ( .A(n1104), .Y(n2422) );
  AND2X1 U1731 ( .A(n2721), .B(DIN[13]), .Y(n1168) );
  INVX1 U1732 ( .A(n1168), .Y(n2423) );
  AND2X1 U1733 ( .A(n2722), .B(DIN[13]), .Y(n1297) );
  INVX1 U1734 ( .A(n1297), .Y(n2424) );
  OR2X1 U1735 ( .A(n1037), .B(n2595), .Y(n2594) );
  OR2X1 U1736 ( .A(n904), .B(n1483), .Y(n2595) );
  AND2X1 U1737 ( .A(n1485), .B(n1306), .Y(n1495) );
  INVX1 U1738 ( .A(n1495), .Y(n2425) );
  AND2X1 U1739 ( .A(n1485), .B(DIN[2]), .Y(n1507) );
  INVX1 U1740 ( .A(n1507), .Y(n2426) );
  AND2X1 U1741 ( .A(n2581), .B(n2132), .Y(n1329) );
  INVX1 U1742 ( .A(n1329), .Y(n2427) );
  AND2X1 U1743 ( .A(n1391), .B(n252), .Y(n1392) );
  INVX1 U1744 ( .A(n1392), .Y(n2428) );
  AND2X1 U1745 ( .A(n1437), .B(n1300), .Y(n1442) );
  INVX1 U1746 ( .A(n1442), .Y(n2429) );
  AND2X1 U1747 ( .A(n1335), .B(DIN[3]), .Y(n1364) );
  INVX1 U1748 ( .A(n1364), .Y(n2430) );
  AND2X1 U1749 ( .A(n2648), .B(n2131), .Y(n1384) );
  INVX1 U1750 ( .A(n1384), .Y(n2431) );
  AND2X1 U1751 ( .A(n2719), .B(n2130), .Y(n1429) );
  INVX1 U1752 ( .A(n1429), .Y(n2432) );
  AND2X1 U1753 ( .A(n2580), .B(n2129), .Y(n1477) );
  INVX1 U1754 ( .A(n1477), .Y(n2433) );
  AND2X1 U1755 ( .A(j_3_), .B(n2666), .Y(n900) );
  INVX1 U1756 ( .A(n900), .Y(n2434) );
  BUFX2 U1757 ( .A(n1194), .Y(n2435) );
  AND2X1 U1758 ( .A(n2647), .B(DIN[14]), .Y(n1105) );
  INVX1 U1759 ( .A(n1105), .Y(n2436) );
  AND2X1 U1760 ( .A(n2711), .B(DIN[13]), .Y(n1075) );
  INVX1 U1761 ( .A(n1075), .Y(n2437) );
  AND2X1 U1762 ( .A(n2710), .B(DIN[13]), .Y(n1139) );
  INVX1 U1763 ( .A(n1139), .Y(n2438) );
  AND2X1 U1764 ( .A(n2650), .B(DIN[15]), .Y(n1233) );
  INVX1 U1765 ( .A(n1233), .Y(n2439) );
  AND2X1 U1766 ( .A(n2649), .B(DIN[14]), .Y(n1298) );
  INVX1 U1767 ( .A(n1298), .Y(n2440) );
  AND2X1 U1768 ( .A(n2712), .B(DIN[13]), .Y(n1268) );
  INVX1 U1769 ( .A(n1268), .Y(n2441) );
  AND2X1 U1770 ( .A(n2655), .B(DIN[10]), .Y(n1277) );
  INVX1 U1771 ( .A(n1277), .Y(n2442) );
  AND2X1 U1772 ( .A(n1142), .B(n1143), .Y(n948) );
  INVX1 U1773 ( .A(n948), .Y(n2443) );
  AND2X1 U1774 ( .A(n1485), .B(DIN[1]), .Y(n1508) );
  INVX1 U1775 ( .A(n1508), .Y(n2444) );
  AND2X1 U1776 ( .A(n2573), .B(n2132), .Y(n1305) );
  INVX1 U1777 ( .A(n1305), .Y(n2445) );
  AND2X1 U1778 ( .A(n2724), .B(n2132), .Y(n1331) );
  INVX1 U1779 ( .A(n1331), .Y(n2446) );
  AND2X1 U1780 ( .A(match_addr[2]), .B(n2827), .Y(n876) );
  INVX1 U1781 ( .A(n876), .Y(n2447) );
  AND2X1 U1782 ( .A(n1391), .B(n1308), .Y(n1403) );
  INVX1 U1783 ( .A(n1403), .Y(n2448) );
  AND2X1 U1784 ( .A(n1437), .B(n252), .Y(n1438) );
  INVX1 U1785 ( .A(n1438), .Y(n2449) );
  AND2X1 U1786 ( .A(n1335), .B(DIN[2]), .Y(n1365) );
  INVX1 U1787 ( .A(n1365), .Y(n2450) );
  AND2X1 U1788 ( .A(n2582), .B(n2131), .Y(n1389) );
  INVX1 U1789 ( .A(n1389), .Y(n2451) );
  AND2X1 U1790 ( .A(n2649), .B(n2130), .Y(n1430) );
  INVX1 U1791 ( .A(n1430), .Y(n2452) );
  AND2X1 U1792 ( .A(n2534), .B(n2129), .Y(n1478) );
  INVX1 U1793 ( .A(n1478), .Y(n2453) );
  AND2X1 U1794 ( .A(n1391), .B(n1306), .Y(n1402) );
  INVX1 U1795 ( .A(n1402), .Y(n2454) );
  AND2X1 U1796 ( .A(n2577), .B(DIN[12]), .Y(n1106) );
  INVX1 U1797 ( .A(n1106), .Y(n2455) );
  AND2X1 U1798 ( .A(n2648), .B(DIN[14]), .Y(n1169) );
  INVX1 U1799 ( .A(n1169), .Y(n2456) );
  AND2X1 U1800 ( .A(n2644), .B(DIN[14]), .Y(n1140) );
  INVX1 U1801 ( .A(n1140), .Y(n2457) );
  AND2X1 U1802 ( .A(n2643), .B(DIN[15]), .Y(n1204) );
  INVX1 U1803 ( .A(n1204), .Y(n2458) );
  AND2X1 U1804 ( .A(n2580), .B(DIN[13]), .Y(n1234) );
  INVX1 U1805 ( .A(n1234), .Y(n2459) );
  AND2X1 U1806 ( .A(n2646), .B(DIN[14]), .Y(n1269) );
  INVX1 U1807 ( .A(n1269), .Y(n2460) );
  AND2X1 U1808 ( .A(n2653), .B(DIN[10]), .Y(n1084) );
  INVX1 U1809 ( .A(n1084), .Y(n2461) );
  AND2X1 U1810 ( .A(n2654), .B(DIN[10]), .Y(n1148) );
  INVX1 U1811 ( .A(n1148), .Y(n2462) );
  AND2X1 U1812 ( .A(n2656), .B(DIN[10]), .Y(n1229) );
  INVX1 U1813 ( .A(n1229), .Y(n2463) );
  AND2X1 U1814 ( .A(n2680), .B(DIN[10]), .Y(n1115) );
  INVX1 U1815 ( .A(n1115), .Y(n2464) );
  AND2X1 U1816 ( .A(n2676), .B(DIN[10]), .Y(n1200) );
  INVX1 U1817 ( .A(n1200), .Y(n2465) );
  AND2X1 U1818 ( .A(n2684), .B(DIN[10]), .Y(n1244) );
  INVX1 U1819 ( .A(n1244), .Y(n2466) );
  AND2X1 U1820 ( .A(n1043), .B(n1044), .Y(n932) );
  INVX1 U1821 ( .A(n932), .Y(n2467) );
  AND2X1 U1822 ( .A(n1271), .B(n1272), .Y(n979) );
  INVX1 U1823 ( .A(n979), .Y(n2468) );
  AND2X1 U1824 ( .A(last[0]), .B(n2848), .Y(n1483) );
  INVX1 U1825 ( .A(n1483), .Y(n2469) );
  BUFX2 U1826 ( .A(n881), .Y(n2470) );
  BUFX2 U1827 ( .A(n988), .Y(n2471) );
  AND2X1 U1828 ( .A(n1485), .B(DIN[0]), .Y(n1509) );
  INVX1 U1829 ( .A(n1509), .Y(n2472) );
  AND2X1 U1830 ( .A(n2716), .B(n2132), .Y(n1317) );
  INVX1 U1831 ( .A(n1317), .Y(n2473) );
  AND2X1 U1832 ( .A(n1391), .B(DIN[4]), .Y(n1412) );
  INVX1 U1833 ( .A(n1412), .Y(n2474) );
  AND2X1 U1834 ( .A(n1437), .B(n1308), .Y(n1449) );
  INVX1 U1835 ( .A(n1449), .Y(n2475) );
  AND2X1 U1836 ( .A(n1335), .B(DIN[1]), .Y(n1366) );
  INVX1 U1837 ( .A(n1366), .Y(n2476) );
  AND2X1 U1838 ( .A(n2725), .B(n2131), .Y(n1390) );
  INVX1 U1839 ( .A(n1390), .Y(n2477) );
  AND2X1 U1840 ( .A(n2575), .B(n2130), .Y(n1423) );
  INVX1 U1841 ( .A(n1423), .Y(n2478) );
  AND2X1 U1842 ( .A(n2655), .B(n2130), .Y(n1434) );
  INVX1 U1843 ( .A(n1434), .Y(n2479) );
  AND2X1 U1844 ( .A(n2584), .B(n2129), .Y(n1481) );
  INVX1 U1845 ( .A(n1481), .Y(n2480) );
  AND2X1 U1846 ( .A(match_addr[1]), .B(n2827), .Y(n873) );
  INVX1 U1847 ( .A(n873), .Y(n2481) );
  AND2X1 U1848 ( .A(n1485), .B(n1302), .Y(n1492) );
  INVX1 U1849 ( .A(n1492), .Y(n2482) );
  AND2X1 U1850 ( .A(n1391), .B(n1304), .Y(n1400) );
  INVX1 U1851 ( .A(n1400), .Y(n2483) );
  AND2X1 U1852 ( .A(n1437), .B(n1306), .Y(n1448) );
  INVX1 U1853 ( .A(n1448), .Y(n2484) );
  AND2X1 U1854 ( .A(n2645), .B(DIN[14]), .Y(n1076) );
  INVX1 U1855 ( .A(n1076), .Y(n2485) );
  AND2X1 U1856 ( .A(n2578), .B(DIN[12]), .Y(n1170) );
  INVX1 U1857 ( .A(n1170), .Y(n2486) );
  AND2X1 U1858 ( .A(n2696), .B(DIN[12]), .Y(n1141) );
  INVX1 U1859 ( .A(n1141), .Y(n2487) );
  AND2X1 U1860 ( .A(n2709), .B(DIN[14]), .Y(n1206) );
  INVX1 U1861 ( .A(n1206), .Y(n2488) );
  AND2X1 U1862 ( .A(n2723), .B(DIN[14]), .Y(n1235) );
  INVX1 U1863 ( .A(n1235), .Y(n2489) );
  AND2X1 U1864 ( .A(n2579), .B(DIN[12]), .Y(n1299) );
  INVX1 U1865 ( .A(n1299), .Y(n2490) );
  AND2X1 U1866 ( .A(n2697), .B(DIN[12]), .Y(n1270) );
  INVX1 U1867 ( .A(n1270), .Y(n2491) );
  AND2X1 U1868 ( .A(n2535), .B(DIN[11]), .Y(n1147) );
  INVX1 U1869 ( .A(n1147), .Y(n2492) );
  AND2X1 U1870 ( .A(n2727), .B(DIN[8]), .Y(n1213) );
  INVX1 U1871 ( .A(n1213), .Y(n2493) );
  AND2X1 U1872 ( .A(n2536), .B(DIN[11]), .Y(n1276) );
  INVX1 U1873 ( .A(n1276), .Y(n2494) );
  AND2X1 U1874 ( .A(n2687), .B(DIN[10]), .Y(n1051) );
  INVX1 U1875 ( .A(n1051), .Y(n2495) );
  AND2X1 U1876 ( .A(n2679), .B(DIN[9]), .Y(n1133) );
  INVX1 U1877 ( .A(n1133), .Y(n2496) );
  AND2X1 U1878 ( .A(n2675), .B(DIN[12]), .Y(n1178) );
  INVX1 U1879 ( .A(n1178), .Y(n2497) );
  AND2X1 U1880 ( .A(n2683), .B(DIN[9]), .Y(n1262) );
  INVX1 U1881 ( .A(n1262), .Y(n2498) );
  BUFX2 U1882 ( .A(n952), .Y(n2499) );
  BUFX2 U1883 ( .A(matchN[0]), .Y(n2500) );
  AND2X1 U1884 ( .A(n1078), .B(n1079), .Y(n914) );
  INVX1 U1885 ( .A(n914), .Y(n2501) );
  AND2X1 U1886 ( .A(n2750), .B(n2585), .Y(n887) );
  INVX1 U1887 ( .A(n887), .Y(n2502) );
  BUFX2 U1888 ( .A(n1522), .Y(n2503) );
  BUFX2 U1889 ( .A(rank[2]), .Y(n2504) );
  AND2X1 U1890 ( .A(n2720), .B(n2132), .Y(n1321) );
  INVX1 U1891 ( .A(n1321), .Y(n2505) );
  AND2X1 U1892 ( .A(n1335), .B(DIN[0]), .Y(n1367) );
  INVX1 U1893 ( .A(n1367), .Y(n2506) );
  AND2X1 U1894 ( .A(n2574), .B(n2131), .Y(n1377) );
  INVX1 U1895 ( .A(n1377), .Y(n2507) );
  AND2X1 U1896 ( .A(n2654), .B(n2131), .Y(n1388) );
  INVX1 U1897 ( .A(n1388), .Y(n2508) );
  AND2X1 U1898 ( .A(n2583), .B(n2130), .Y(n1435) );
  INVX1 U1899 ( .A(n1435), .Y(n2509) );
  AND2X1 U1900 ( .A(n2576), .B(n2129), .Y(n1468) );
  INVX1 U1901 ( .A(n1468), .Y(n2510) );
  AND2X1 U1902 ( .A(n2718), .B(n2129), .Y(n1479) );
  INVX1 U1903 ( .A(n1479), .Y(n2511) );
  AND2X1 U1904 ( .A(match_addr[0]), .B(n2827), .Y(n870) );
  INVX1 U1905 ( .A(n870), .Y(n2512) );
  AND2X1 U1906 ( .A(n1485), .B(n1300), .Y(n1490) );
  INVX1 U1907 ( .A(n1490), .Y(n2513) );
  AND2X1 U1908 ( .A(n1391), .B(n250), .Y(n1395) );
  INVX1 U1909 ( .A(n1395), .Y(n2514) );
  AND2X1 U1910 ( .A(n1437), .B(DIN[6]), .Y(n1455) );
  INVX1 U1911 ( .A(n1455), .Y(n2515) );
  AND2X1 U1912 ( .A(n1437), .B(n1304), .Y(n1446) );
  INVX1 U1913 ( .A(n1446), .Y(n2516) );
  AND2X1 U1914 ( .A(n1335), .B(n1302), .Y(n1342) );
  INVX1 U1915 ( .A(n1342), .Y(n2517) );
  AND2X1 U1916 ( .A(n2698), .B(DIN[12]), .Y(n1077) );
  INVX1 U1917 ( .A(n1077), .Y(n2518) );
  AND2X1 U1918 ( .A(n2695), .B(DIN[13]), .Y(n1205) );
  INVX1 U1919 ( .A(n1205), .Y(n2519) );
  AND2X1 U1920 ( .A(n2724), .B(DIN[8]), .Y(n1100) );
  INVX1 U1921 ( .A(n1100), .Y(n2520) );
  AND2X1 U1922 ( .A(n2725), .B(DIN[8]), .Y(n1164) );
  INVX1 U1923 ( .A(n1164), .Y(n2521) );
  AND2X1 U1924 ( .A(n2726), .B(DIN[8]), .Y(n1293) );
  INVX1 U1925 ( .A(n1293), .Y(n2522) );
  AND2X1 U1926 ( .A(n2584), .B(DIN[9]), .Y(n1228) );
  INVX1 U1927 ( .A(n1228), .Y(n2523) );
  AND2X1 U1928 ( .A(n2688), .B(DIN[9]), .Y(n1069) );
  INVX1 U1929 ( .A(n1069), .Y(n2524) );
  BUFX2 U1930 ( .A(n983), .Y(n2525) );
  AND2X1 U1931 ( .A(n1107), .B(n1108), .Y(n964) );
  INVX1 U1932 ( .A(n964), .Y(n2526) );
  AND2X1 U1933 ( .A(n1236), .B(n1237), .Y(n995) );
  INVX1 U1934 ( .A(n995), .Y(n2527) );
  OR2X1 U1935 ( .A(n2800), .B(n2798), .Y(n885) );
  INVX1 U1936 ( .A(n885), .Y(n2528) );
  BUFX2 U1937 ( .A(mem[126]), .Y(n2529) );
  BUFX2 U1938 ( .A(mem[94]), .Y(n2530) );
  BUFX2 U1939 ( .A(mem[62]), .Y(n2531) );
  BUFX2 U1940 ( .A(mem[31]), .Y(n2532) );
  BUFX2 U1941 ( .A(mem[115]), .Y(n2533) );
  BUFX2 U1942 ( .A(mem[20]), .Y(n2534) );
  BUFX2 U1943 ( .A(mem[83]), .Y(n2535) );
  BUFX2 U1944 ( .A(mem[51]), .Y(n2536) );
  INVX1 U1945 ( .A(n1003), .Y(n2537) );
  BUFX2 U1946 ( .A(n1018), .Y(n2538) );
  BUFX2 U1947 ( .A(matchN[4]), .Y(n2539) );
  BUFX2 U1948 ( .A(n1513), .Y(n2540) );
  BUFX2 U1949 ( .A(rank[20]), .Y(n2541) );
  BUFX2 U1950 ( .A(rank[17]), .Y(n2542) );
  BUFX2 U1951 ( .A(rank[1]), .Y(n2543) );
  BUFX2 U1952 ( .A(n1334), .Y(n2544) );
  AND2X1 U1953 ( .A(n2647), .B(n2132), .Y(n1319) );
  INVX1 U1954 ( .A(n1319), .Y(n2545) );
  AND2X1 U1955 ( .A(n2721), .B(n2131), .Y(n1385) );
  INVX1 U1956 ( .A(n1385), .Y(n2546) );
  AND2X1 U1957 ( .A(n2726), .B(n2130), .Y(n1436) );
  INVX1 U1958 ( .A(n1436), .Y(n2547) );
  AND2X1 U1959 ( .A(n2642), .B(n2129), .Y(n1469) );
  INVX1 U1960 ( .A(n1469), .Y(n2548) );
  AND2X1 U1961 ( .A(n2656), .B(n2129), .Y(n1480) );
  INVX1 U1962 ( .A(n1480), .Y(n2549) );
  AND2X1 U1963 ( .A(n1485), .B(DIN[7]), .Y(n1501) );
  INVX1 U1964 ( .A(n1501), .Y(n2550) );
  AND2X1 U1965 ( .A(n1391), .B(DIN[6]), .Y(n1409) );
  INVX1 U1966 ( .A(n1409), .Y(n2551) );
  AND2X1 U1967 ( .A(n1391), .B(n1302), .Y(n1398) );
  INVX1 U1968 ( .A(n1398), .Y(n2552) );
  AND2X1 U1969 ( .A(n1437), .B(n250), .Y(n1441) );
  INVX1 U1970 ( .A(n1441), .Y(n2553) );
  AND2X1 U1971 ( .A(n1335), .B(n1304), .Y(n1345) );
  INVX1 U1972 ( .A(n1345), .Y(n2554) );
  AND2X1 U1973 ( .A(n1335), .B(DIN[6]), .Y(n1360) );
  INVX1 U1974 ( .A(n1360), .Y(n2555) );
  INVX1 U1975 ( .A(n1781), .Y(n2556) );
  INVX1 U1976 ( .A(n874), .Y(n2557) );
  INVX1 U1977 ( .A(n2984), .Y(n2558) );
  AND2X1 U1978 ( .A(n2699), .B(n2622), .Y(n2984) );
  INVX1 U1979 ( .A(n1083), .Y(n2559) );
  AND2X1 U1980 ( .A(n2689), .B(DIN[8]), .Y(n1071) );
  INVX1 U1981 ( .A(n1071), .Y(n2560) );
  AND2X1 U1982 ( .A(n2678), .B(DIN[8]), .Y(n1135) );
  INVX1 U1983 ( .A(n1135), .Y(n2561) );
  AND2X1 U1984 ( .A(n2677), .B(DIN[8]), .Y(n1180) );
  INVX1 U1985 ( .A(n1180), .Y(n2562) );
  AND2X1 U1986 ( .A(n2682), .B(DIN[8]), .Y(n1264) );
  INVX1 U1987 ( .A(n1264), .Y(n2563) );
  AND2X1 U1988 ( .A(n2657), .B(n2774), .Y(n1648) );
  INVX1 U1989 ( .A(n1648), .Y(n2564) );
  BUFX2 U1990 ( .A(mem[122]), .Y(n2565) );
  BUFX2 U1991 ( .A(mem[90]), .Y(n2566) );
  BUFX2 U1992 ( .A(mem[58]), .Y(n2567) );
  BUFX2 U1993 ( .A(mem[26]), .Y(n2568) );
  BUFX2 U1994 ( .A(mem[15]), .Y(n2569) );
  BUFX2 U1995 ( .A(mem[76]), .Y(n2570) );
  BUFX2 U1996 ( .A(mem[44]), .Y(n2571) );
  BUFX2 U1997 ( .A(mem[110]), .Y(n2572) );
  BUFX2 U1998 ( .A(mem[125]), .Y(n2573) );
  BUFX2 U1999 ( .A(mem[93]), .Y(n2574) );
  BUFX2 U2000 ( .A(mem[61]), .Y(n2575) );
  BUFX2 U2001 ( .A(mem[30]), .Y(n2576) );
  BUFX2 U2002 ( .A(mem[116]), .Y(n2577) );
  BUFX2 U2003 ( .A(mem[84]), .Y(n2578) );
  BUFX2 U2004 ( .A(mem[52]), .Y(n2579) );
  BUFX2 U2005 ( .A(mem[21]), .Y(n2580) );
  BUFX2 U2006 ( .A(mem[113]), .Y(n2581) );
  BUFX2 U2007 ( .A(mem[81]), .Y(n2582) );
  BUFX2 U2008 ( .A(mem[49]), .Y(n2583) );
  BUFX2 U2009 ( .A(mem[17]), .Y(n2584) );
  BUFX2 U2010 ( .A(n906), .Y(n2585) );
  AND2X1 U2011 ( .A(n2809), .B(n967), .Y(n976) );
  INVX1 U2012 ( .A(n976), .Y(n2586) );
  BUFX2 U2013 ( .A(rank[23]), .Y(n2587) );
  BUFX2 U2014 ( .A(rank[14]), .Y(n2588) );
  BUFX2 U2015 ( .A(rank[5]), .Y(n2589) );
  BUFX2 U2016 ( .A(rank[11]), .Y(n2590) );
  BUFX2 U2017 ( .A(n1005), .Y(n2591) );
  AND2X1 U2018 ( .A(n998), .B(n2961), .Y(n1009) );
  INVX1 U2019 ( .A(n1009), .Y(n2592) );
  AND2X1 U2020 ( .A(n2674), .B(n1003), .Y(n998) );
  BUFX2 U2021 ( .A(rank[7]), .Y(n2593) );
  BUFX2 U2022 ( .A(rank[0]), .Y(n2596) );
  BUFX2 U2023 ( .A(n886), .Y(n2597) );
  AND2X1 U2024 ( .A(n2805), .B(n936), .Y(n945) );
  INVX1 U2025 ( .A(n945), .Y(n2598) );
  AND2X1 U2026 ( .A(n2700), .B(n2132), .Y(n1027) );
  INVX1 U2027 ( .A(n1027), .Y(n2599) );
  AND2X1 U2028 ( .A(n2717), .B(n2131), .Y(n1383) );
  INVX1 U2029 ( .A(n1383), .Y(n2600) );
  AND2X1 U2030 ( .A(n2722), .B(n2130), .Y(n1431) );
  INVX1 U2031 ( .A(n1431), .Y(n2601) );
  AND2X1 U2032 ( .A(n2727), .B(n2129), .Y(n1482) );
  INVX1 U2033 ( .A(n1482), .Y(n2602) );
  AND2X1 U2034 ( .A(n1485), .B(n1304), .Y(n1494) );
  INVX1 U2035 ( .A(n1494), .Y(n2603) );
  AND2X1 U2036 ( .A(n1485), .B(DIN[6]), .Y(n1503) );
  INVX1 U2037 ( .A(n1503), .Y(n2604) );
  AND2X1 U2038 ( .A(n1391), .B(DIN[5]), .Y(n1411) );
  INVX1 U2039 ( .A(n1411), .Y(n2605) );
  AND2X1 U2040 ( .A(n1437), .B(DIN[5]), .Y(n1457) );
  INVX1 U2041 ( .A(n1457), .Y(n2606) );
  AND2X1 U2042 ( .A(n1437), .B(n1302), .Y(n1444) );
  INVX1 U2043 ( .A(n1444), .Y(n2607) );
  AND2X1 U2044 ( .A(n1335), .B(n1306), .Y(n1348) );
  INVX1 U2045 ( .A(n1348), .Y(n2608) );
  AND2X1 U2046 ( .A(n1335), .B(DIN[5]), .Y(n1362) );
  INVX1 U2047 ( .A(n1362), .Y(n2609) );
  BUFX2 U2048 ( .A(n3000), .Y(match_addr[2]) );
  BUFX2 U2049 ( .A(n3001), .Y(match_addr[1]) );
  BUFX2 U2050 ( .A(n3002), .Y(match_addr[0]) );
  AND2X1 U2051 ( .A(n2686), .B(DIN[11]), .Y(n1049) );
  INVX1 U2052 ( .A(n1049), .Y(n2613) );
  AND2X1 U2053 ( .A(n2681), .B(DIN[11]), .Y(n1113) );
  INVX1 U2054 ( .A(n1113), .Y(n2614) );
  AND2X1 U2055 ( .A(n2685), .B(DIN[11]), .Y(n1242) );
  INVX1 U2056 ( .A(n1242), .Y(n2615) );
  AND2X1 U2057 ( .A(n2692), .B(DIN[9]), .Y(n1198) );
  INVX1 U2058 ( .A(n1198), .Y(n2616) );
  BUFX2 U2059 ( .A(m), .Y(n2617) );
  BUFX2 U2060 ( .A(mem[127]), .Y(n2618) );
  BUFX2 U2061 ( .A(mem[95]), .Y(n2619) );
  BUFX2 U2062 ( .A(mem[27]), .Y(n2620) );
  BUFX2 U2063 ( .A(mem[63]), .Y(n2621) );
  AND2X1 U2064 ( .A(n236), .B(n2823), .Y(n2986) );
  INVX1 U2065 ( .A(n2986), .Y(n2622) );
  BUFX2 U2066 ( .A(mem[123]), .Y(n2623) );
  BUFX2 U2067 ( .A(mem[91]), .Y(n2624) );
  BUFX2 U2068 ( .A(mem[59]), .Y(n2625) );
  BUFX2 U2069 ( .A(mem[121]), .Y(n2626) );
  BUFX2 U2070 ( .A(mem[120]), .Y(n2627) );
  BUFX2 U2071 ( .A(mem[89]), .Y(n2628) );
  BUFX2 U2072 ( .A(mem[88]), .Y(n2629) );
  BUFX2 U2073 ( .A(mem[57]), .Y(n2630) );
  BUFX2 U2074 ( .A(mem[56]), .Y(n2631) );
  BUFX2 U2075 ( .A(mem[28]), .Y(n2632) );
  BUFX2 U2076 ( .A(mem[24]), .Y(n2633) );
  BUFX2 U2077 ( .A(mem[25]), .Y(n2634) );
  BUFX2 U2078 ( .A(mem[14]), .Y(n2635) );
  BUFX2 U2079 ( .A(mem[77]), .Y(n2636) );
  BUFX2 U2080 ( .A(mem[45]), .Y(n2637) );
  BUFX2 U2081 ( .A(mem[109]), .Y(n2638) );
  BUFX2 U2082 ( .A(mem[124]), .Y(n2639) );
  BUFX2 U2083 ( .A(mem[92]), .Y(n2640) );
  BUFX2 U2084 ( .A(mem[60]), .Y(n2641) );
  BUFX2 U2085 ( .A(mem[29]), .Y(n2642) );
  BUFX2 U2086 ( .A(mem[7]), .Y(n2643) );
  BUFX2 U2087 ( .A(mem[70]), .Y(n2644) );
  BUFX2 U2088 ( .A(mem[102]), .Y(n2645) );
  BUFX2 U2089 ( .A(mem[38]), .Y(n2646) );
  BUFX2 U2090 ( .A(mem[118]), .Y(n2647) );
  BUFX2 U2091 ( .A(mem[86]), .Y(n2648) );
  BUFX2 U2092 ( .A(mem[54]), .Y(n2649) );
  BUFX2 U2093 ( .A(mem[23]), .Y(n2650) );
  BUFX2 U2094 ( .A(matchN[12]), .Y(n2651) );
  BUFX2 U2095 ( .A(matchN[6]), .Y(n2652) );
  BUFX2 U2096 ( .A(mem[114]), .Y(n2653) );
  BUFX2 U2097 ( .A(mem[82]), .Y(n2654) );
  BUFX2 U2098 ( .A(mem[50]), .Y(n2655) );
  BUFX2 U2099 ( .A(mem[18]), .Y(n2656) );
  BUFX2 U2100 ( .A(rank[8]), .Y(n2657) );
  BUFX2 U2101 ( .A(rank[22]), .Y(n2658) );
  BUFX2 U2102 ( .A(rank[13]), .Y(n2659) );
  BUFX2 U2103 ( .A(rank[4]), .Y(n2660) );
  BUFX2 U2104 ( .A(rank[10]), .Y(n2661) );
  BUFX2 U2105 ( .A(matchN[3]), .Y(n2662) );
  BUFX2 U2106 ( .A(rank[18]), .Y(n2663) );
  BUFX2 U2107 ( .A(rank[15]), .Y(n2664) );
  BUFX2 U2108 ( .A(n1369), .Y(n2665) );
  AND2X1 U2109 ( .A(n2793), .B(n901), .Y(n880) );
  INVX1 U2110 ( .A(n880), .Y(n2666) );
  INVX1 U2111 ( .A(n905), .Y(n2667) );
  AND2X1 U2112 ( .A(n1437), .B(n251), .Y(n1439) );
  INVX1 U2113 ( .A(n1439), .Y(n2668) );
  AND2X1 U2114 ( .A(n1335), .B(n250), .Y(n1338) );
  INVX1 U2115 ( .A(n1338), .Y(n2669) );
  INVX1 U2116 ( .A(n1099), .Y(n2670) );
  INVX1 U2117 ( .A(n1163), .Y(n2671) );
  INVX1 U2118 ( .A(n1212), .Y(n2672) );
  INVX1 U2119 ( .A(n1292), .Y(n2673) );
  BUFX2 U2120 ( .A(matchN[2]), .Y(n2674) );
  BUFX2 U2121 ( .A(mem[4]), .Y(n2675) );
  BUFX2 U2122 ( .A(mem[2]), .Y(n2676) );
  BUFX2 U2123 ( .A(mem[0]), .Y(n2677) );
  BUFX2 U2124 ( .A(mem[64]), .Y(n2678) );
  BUFX2 U2125 ( .A(mem[65]), .Y(n2679) );
  BUFX2 U2126 ( .A(mem[66]), .Y(n2680) );
  BUFX2 U2127 ( .A(mem[67]), .Y(n2681) );
  BUFX2 U2128 ( .A(mem[32]), .Y(n2682) );
  BUFX2 U2129 ( .A(mem[33]), .Y(n2683) );
  BUFX2 U2130 ( .A(mem[34]), .Y(n2684) );
  BUFX2 U2131 ( .A(mem[35]), .Y(n2685) );
  BUFX2 U2132 ( .A(mem[99]), .Y(n2686) );
  BUFX2 U2133 ( .A(mem[98]), .Y(n2687) );
  BUFX2 U2134 ( .A(mem[97]), .Y(n2688) );
  BUFX2 U2135 ( .A(mem[96]), .Y(n2689) );
  BUFX2 U2136 ( .A(matchN[16]), .Y(n2690) );
  BUFX2 U2137 ( .A(matchN[10]), .Y(n2691) );
  BUFX2 U2138 ( .A(mem[1]), .Y(n2692) );
  BUFX2 U2139 ( .A(matchN[23]), .Y(n2693) );
  BUFX2 U2140 ( .A(matchN[22]), .Y(n2694) );
  BUFX2 U2141 ( .A(mem[5]), .Y(n2695) );
  BUFX2 U2142 ( .A(mem[68]), .Y(n2696) );
  BUFX2 U2143 ( .A(mem[36]), .Y(n2697) );
  BUFX2 U2144 ( .A(mem[100]), .Y(n2698) );
  AND2X1 U2145 ( .A(n2987), .B(n2988), .Y(n2985) );
  INVX1 U2146 ( .A(n2985), .Y(n2699) );
  BUFX2 U2147 ( .A(matchN[21]), .Y(n2700) );
  BUFX2 U2148 ( .A(mem[3]), .Y(n2701) );
  BUFX2 U2149 ( .A(mem[71]), .Y(n2702) );
  BUFX2 U2150 ( .A(mem[103]), .Y(n2703) );
  BUFX2 U2151 ( .A(mem[39]), .Y(n2704) );
  BUFX2 U2152 ( .A(mem[13]), .Y(n2705) );
  BUFX2 U2153 ( .A(mem[78]), .Y(n2706) );
  BUFX2 U2154 ( .A(mem[46]), .Y(n2707) );
  BUFX2 U2155 ( .A(mem[108]), .Y(n2708) );
  BUFX2 U2156 ( .A(mem[6]), .Y(n2709) );
  BUFX2 U2157 ( .A(mem[69]), .Y(n2710) );
  BUFX2 U2158 ( .A(mem[101]), .Y(n2711) );
  BUFX2 U2159 ( .A(mem[37]), .Y(n2712) );
  BUFX2 U2160 ( .A(matchN[17]), .Y(n2713) );
  BUFX2 U2161 ( .A(matchN[11]), .Y(n2714) );
  BUFX2 U2162 ( .A(matchN[5]), .Y(n2715) );
  BUFX2 U2163 ( .A(mem[119]), .Y(n2716) );
  BUFX2 U2164 ( .A(mem[87]), .Y(n2717) );
  BUFX2 U2165 ( .A(mem[19]), .Y(n2718) );
  BUFX2 U2166 ( .A(mem[55]), .Y(n2719) );
  BUFX2 U2167 ( .A(mem[117]), .Y(n2720) );
  BUFX2 U2168 ( .A(mem[85]), .Y(n2721) );
  BUFX2 U2169 ( .A(mem[53]), .Y(n2722) );
  BUFX2 U2170 ( .A(mem[22]), .Y(n2723) );
  BUFX2 U2171 ( .A(mem[112]), .Y(n2724) );
  BUFX2 U2172 ( .A(mem[80]), .Y(n2725) );
  BUFX2 U2173 ( .A(mem[48]), .Y(n2726) );
  BUFX2 U2174 ( .A(mem[16]), .Y(n2727) );
  BUFX2 U2175 ( .A(matchN[15]), .Y(n2728) );
  BUFX2 U2176 ( .A(matchN[9]), .Y(n2729) );
  AND2X1 U2177 ( .A(EN), .B(n2946), .Y(n903) );
  INVX1 U2178 ( .A(n903), .Y(n2730) );
  BUFX2 U2179 ( .A(rank[19]), .Y(n2731) );
  BUFX2 U2180 ( .A(rank[16]), .Y(n2732) );
  BUFX2 U2181 ( .A(matchN[1]), .Y(n2733) );
  BUFX2 U2182 ( .A(rank[21]), .Y(n2734) );
  BUFX2 U2183 ( .A(rank[12]), .Y(n2735) );
  BUFX2 U2184 ( .A(rank[3]), .Y(n2736) );
  BUFX2 U2185 ( .A(rank[6]), .Y(n2737) );
  BUFX2 U2186 ( .A(rank[9]), .Y(n2738) );
  AND2X1 U2187 ( .A(DIN[3]), .B(DIN[11]), .Y(n1308) );
  INVX1 U2188 ( .A(n1308), .Y(n2739) );
  AND2X1 U2189 ( .A(DIN[2]), .B(DIN[10]), .Y(n1310) );
  INVX1 U2190 ( .A(n1310), .Y(n2740) );
  AND2X1 U2191 ( .A(DIN[1]), .B(DIN[9]), .Y(n1312) );
  INVX1 U2192 ( .A(n1312), .Y(n2741) );
  AND2X1 U2193 ( .A(DIN[0]), .B(DIN[8]), .Y(n1314) );
  INVX1 U2194 ( .A(n1314), .Y(n2742) );
  AND2X1 U2195 ( .A(DIN[7]), .B(DIN[15]), .Y(n1300) );
  INVX1 U2196 ( .A(n1300), .Y(n2743) );
  AND2X1 U2197 ( .A(DIN[4]), .B(DIN[12]), .Y(n1306) );
  INVX1 U2198 ( .A(n1306), .Y(n2744) );
  AND2X1 U2199 ( .A(DIN[6]), .B(DIN[14]), .Y(n1302) );
  INVX1 U2200 ( .A(n1302), .Y(n2745) );
  AND2X1 U2201 ( .A(DIN[5]), .B(DIN[13]), .Y(n1304) );
  INVX1 U2202 ( .A(n1304), .Y(n2746) );
  BUFX2 U2203 ( .A(n1368), .Y(n2747) );
  BUFX2 U2204 ( .A(n892), .Y(n2748) );
  AND2X1 U2205 ( .A(n2803), .B(n2802), .Y(n929) );
  INVX1 U2206 ( .A(n929), .Y(n2749) );
  BUFX2 U2207 ( .A(n897), .Y(n2750) );
  AND2X1 U2208 ( .A(n2810), .B(n2811), .Y(n992) );
  INVX1 U2209 ( .A(n992), .Y(n2751) );
  INVX1 U2210 ( .A(n868), .Y(n2752) );
  BUFX2 U2211 ( .A(n888), .Y(n2753) );
  AND2X1 U2212 ( .A(n2807), .B(n2806), .Y(n961) );
  INVX1 U2213 ( .A(n961), .Y(n2754) );
  INVX1 U2214 ( .A(n251), .Y(n2813) );
  INVX1 U2215 ( .A(n252), .Y(n2814) );
  INVX1 U2216 ( .A(n2794), .Y(n2793) );
  INVX1 U2217 ( .A(n2794), .Y(n2792) );
  INVX1 U2218 ( .A(n2794), .Y(n2791) );
  INVX1 U2219 ( .A(reset), .Y(n2790) );
  INVX1 U2220 ( .A(reset), .Y(n2789) );
  INVX1 U2221 ( .A(reset), .Y(n2788) );
  INVX1 U2222 ( .A(reset), .Y(n2787) );
  INVX1 U2223 ( .A(reset), .Y(n2785) );
  INVX1 U2224 ( .A(reset), .Y(n2786) );
  INVX1 U2225 ( .A(reset), .Y(n2784) );
  INVX1 U2226 ( .A(reset), .Y(n2783) );
  INVX1 U2227 ( .A(reset), .Y(n2782) );
  INVX1 U2228 ( .A(reset), .Y(n2781) );
  INVX1 U2229 ( .A(reset), .Y(n2780) );
  INVX1 U2230 ( .A(reset), .Y(n2779) );
  INVX1 U2231 ( .A(n2597), .Y(n2804) );
  INVX1 U2232 ( .A(n2748), .Y(n2800) );
  INVX1 U2233 ( .A(n2585), .Y(n2808) );
  INVX1 U2234 ( .A(n2753), .Y(n2801) );
  INVX1 U2235 ( .A(n250), .Y(n2816) );
  INVX1 U2236 ( .A(n1660), .Y(n2832) );
  INVX1 U2237 ( .A(n1617), .Y(n2836) );
  INVX1 U2238 ( .A(n1639), .Y(n2834) );
  INVX1 U2239 ( .A(n1596), .Y(n2838) );
  INVX1 U2240 ( .A(n1534), .Y(n2830) );
  INVX1 U2241 ( .A(n1575), .Y(n2840) );
  INVX1 U2242 ( .A(n1548), .Y(n2842) );
  INVX1 U2243 ( .A(n1681), .Y(n2828) );
  BUFX2 U2244 ( .A(n904), .Y(n2775) );
  BUFX2 U2245 ( .A(n904), .Y(n2776) );
  INVX1 U2246 ( .A(n2777), .Y(n2794) );
  INVX1 U2247 ( .A(n1037), .Y(n2873) );
  INVX1 U2248 ( .A(n2591), .Y(n2812) );
  OR2X1 U2249 ( .A(n2878), .B(n912), .Y(n916) );
  INVX1 U2250 ( .A(n2306), .Y(n2802) );
  INVX1 U2251 ( .A(n2499), .Y(n2806) );
  INVX1 U2252 ( .A(n2525), .Y(n2811) );
  INVX1 U2253 ( .A(n2133), .Y(n2798) );
  AND2X1 U2254 ( .A(n1172), .B(n1173), .Y(n1017) );
  AND2X1 U2255 ( .A(n235), .B(n233), .Y(n2987) );
  INVX1 U2256 ( .A(n2778), .Y(n2777) );
  INVX1 U2257 ( .A(n2503), .Y(n2874) );
  INVX1 U2258 ( .A(n2747), .Y(n2846) );
  INVX1 U2259 ( .A(n2665), .Y(n2847) );
  INVX1 U2260 ( .A(n2715), .Y(n2961) );
  INVX1 U2261 ( .A(n2539), .Y(n2962) );
  INVX1 U2262 ( .A(n2718), .Y(n2966) );
  AND2X1 U2263 ( .A(DIN[11]), .B(n2859), .Y(n1183) );
  INVX1 U2264 ( .A(n953), .Y(n2805) );
  INVX1 U2265 ( .A(n2470), .Y(n2797) );
  INVX1 U2266 ( .A(n984), .Y(n2809) );
  OR2X1 U2267 ( .A(n2879), .B(n919), .Y(n917) );
  INVX1 U2268 ( .A(n2074), .Y(n2799) );
  INVX1 U2269 ( .A(n999), .Y(n2810) );
  INVX1 U2270 ( .A(n968), .Y(n2807) );
  INVX1 U2271 ( .A(n937), .Y(n2803) );
  AND2X1 U2272 ( .A(n1207), .B(n1208), .Y(n1011) );
  AND2X1 U2273 ( .A(DIN[11]), .B(n2963), .Y(n1216) );
  INVX1 U2274 ( .A(n2134), .Y(n2795) );
  AND2X1 U2275 ( .A(DIN[15]), .B(n2924), .Y(n1247) );
  INVX1 U2276 ( .A(n2719), .Y(n2957) );
  INVX1 U2277 ( .A(n2717), .Y(n2950) );
  AND2X1 U2278 ( .A(DIN[15]), .B(n2905), .Y(n1118) );
  INVX1 U2279 ( .A(n2580), .Y(n2964) );
  INVX1 U2280 ( .A(n2534), .Y(n2965) );
  INVX1 U2281 ( .A(n2733), .Y(n2853) );
  INVX1 U2282 ( .A(n2500), .Y(n2854) );
  INVX1 U2283 ( .A(n1221), .Y(n2967) );
  INVX1 U2284 ( .A(n2084), .Y(n2924) );
  INVX1 U2285 ( .A(n2099), .Y(n2859) );
  INVX1 U2286 ( .A(n2701), .Y(n2867) );
  INVX1 U2287 ( .A(n2620), .Y(n2963) );
  INVX1 U2288 ( .A(n2682), .Y(n2909) );
  INVX1 U2289 ( .A(n2677), .Y(n2870) );
  INVX1 U2290 ( .A(n2697), .Y(n2913) );
  INVX1 U2291 ( .A(n2684), .Y(n2911) );
  INVX1 U2292 ( .A(n2695), .Y(n2865) );
  INVX1 U2293 ( .A(n2676), .Y(n2868) );
  INVX1 U2294 ( .A(n2685), .Y(n2912) );
  INVX1 U2295 ( .A(n2683), .Y(n2910) );
  INVX1 U2296 ( .A(n2675), .Y(n2866) );
  INVX1 U2297 ( .A(n2692), .Y(n2869) );
  INVX1 U2298 ( .A(n2674), .Y(n2852) );
  INVX1 U2299 ( .A(n2096), .Y(n2862) );
  INVX1 U2300 ( .A(n2100), .Y(n2858) );
  INVX1 U2301 ( .A(n2098), .Y(n2860) );
  INVX1 U2302 ( .A(n2097), .Y(n2861) );
  AND2X1 U2303 ( .A(DIN[15]), .B(n2956), .Y(n1280) );
  AND2X1 U2304 ( .A(DIN[15]), .B(n2949), .Y(n1151) );
  AND2X1 U2305 ( .A(DIN[15]), .B(n2930), .Y(n1054) );
  INVX1 U2306 ( .A(n2716), .Y(n2881) );
  INVX1 U2307 ( .A(n2709), .Y(n2864) );
  INVX1 U2308 ( .A(n2643), .Y(n2863) );
  INVX1 U2309 ( .A(n2705), .Y(n2857) );
  INVX1 U2310 ( .A(n2635), .Y(n2856) );
  INVX1 U2311 ( .A(n2569), .Y(n2855) );
  INVX1 U2312 ( .A(n2646), .Y(n2915) );
  INVX1 U2313 ( .A(n2712), .Y(n2914) );
  INVX1 U2314 ( .A(n2644), .Y(n2896) );
  INVX1 U2315 ( .A(n2710), .Y(n2895) );
  INVX1 U2316 ( .A(n2711), .Y(n2940) );
  INVX1 U2317 ( .A(n2645), .Y(n2939) );
  INVX1 U2318 ( .A(n2652), .Y(n2925) );
  INVX1 U2319 ( .A(n2707), .Y(n2923) );
  INVX1 U2320 ( .A(n2637), .Y(n2922) );
  INVX1 U2321 ( .A(n2571), .Y(n2921) );
  INVX1 U2322 ( .A(n2651), .Y(n2906) );
  INVX1 U2323 ( .A(n2706), .Y(n2904) );
  INVX1 U2324 ( .A(n2636), .Y(n2903) );
  INVX1 U2325 ( .A(n2570), .Y(n2902) );
  INVX1 U2326 ( .A(n2708), .Y(n2933) );
  INVX1 U2327 ( .A(n2638), .Y(n2932) );
  INVX1 U2328 ( .A(n2572), .Y(n2931) );
  INVX1 U2329 ( .A(n1657), .Y(n2833) );
  INVX1 U2330 ( .A(n1614), .Y(n2837) );
  INVX1 U2331 ( .A(n1636), .Y(n2835) );
  INVX1 U2332 ( .A(n1593), .Y(n2839) );
  INVX1 U2333 ( .A(n1533), .Y(n2831) );
  INVX1 U2334 ( .A(n1572), .Y(n2841) );
  INVX1 U2335 ( .A(n1545), .Y(n2843) );
  INVX1 U2336 ( .A(n1678), .Y(n2829) );
  INVX1 U2337 ( .A(n2579), .Y(n2958) );
  INVX1 U2338 ( .A(n2536), .Y(n2959) );
  INVX1 U2339 ( .A(n2578), .Y(n2951) );
  INVX1 U2340 ( .A(n2535), .Y(n2952) );
  INVX1 U2341 ( .A(last[1]), .Y(n2889) );
  INVX1 U2342 ( .A(last[2]), .Y(n2877) );
  INVX1 U2343 ( .A(last[0]), .Y(n2851) );
  INVX1 U2344 ( .A(n1285), .Y(n2960) );
  INVX1 U2345 ( .A(n1156), .Y(n2953) );
  INVX1 U2346 ( .A(n2083), .Y(n2926) );
  INVX1 U2347 ( .A(n2090), .Y(n2907) );
  INVX1 U2348 ( .A(n2101), .Y(n2815) );
  AND2X1 U2349 ( .A(DIN[4]), .B(n238), .Y(n2992) );
  INVX1 U2350 ( .A(n2102), .Y(n2818) );
  AND2X1 U2351 ( .A(DIN[6]), .B(DIN[5]), .Y(n2995) );
  INVX1 U2352 ( .A(n2103), .Y(n2823) );
  AND2X1 U2353 ( .A(DIN[1]), .B(DIN[2]), .Y(n2998) );
  INVX1 U2354 ( .A(n2691), .Y(n2955) );
  INVX1 U2355 ( .A(n2690), .Y(n2948) );
  INVX1 U2356 ( .A(n2091), .Y(n2905) );
  INVX1 U2357 ( .A(n2704), .Y(n2916) );
  INVX1 U2358 ( .A(n2702), .Y(n2897) );
  INVX1 U2359 ( .A(n2714), .Y(n2954) );
  INVX1 U2360 ( .A(n2713), .Y(n2947) );
  INVX1 U2361 ( .A(n2621), .Y(n2956) );
  INVX1 U2362 ( .A(n2619), .Y(n2949) );
  INVX1 U2363 ( .A(n2678), .Y(n2890) );
  INVX1 U2364 ( .A(n2696), .Y(n2894) );
  INVX1 U2365 ( .A(n2680), .Y(n2892) );
  INVX1 U2366 ( .A(n2681), .Y(n2893) );
  INVX1 U2367 ( .A(n2679), .Y(n2891) );
  INVX1 U2368 ( .A(DIN[0]), .Y(n2826) );
  INVX1 U2369 ( .A(DIN[1]), .Y(n2825) );
  INVX1 U2370 ( .A(DIN[2]), .Y(n2824) );
  INVX1 U2371 ( .A(DIN[3]), .Y(n2822) );
  INVX1 U2372 ( .A(DIN[4]), .Y(n2821) );
  INVX1 U2373 ( .A(DIN[5]), .Y(n2820) );
  INVX1 U2374 ( .A(DIN[6]), .Y(n2819) );
  INVX1 U2375 ( .A(DIN[7]), .Y(n2817) );
  INVX1 U2376 ( .A(n2088), .Y(n2917) );
  INVX1 U2377 ( .A(n2087), .Y(n2918) );
  INVX1 U2378 ( .A(n2086), .Y(n2919) );
  INVX1 U2379 ( .A(n2085), .Y(n2920) );
  INVX1 U2380 ( .A(n2095), .Y(n2898) );
  INVX1 U2381 ( .A(n2094), .Y(n2899) );
  INVX1 U2382 ( .A(n2093), .Y(n2900) );
  INVX1 U2383 ( .A(n2092), .Y(n2901) );
  INVX1 U2384 ( .A(n2082), .Y(n2927) );
  INVX1 U2385 ( .A(n2089), .Y(n2908) );
  AND2X1 U2386 ( .A(DIN[15]), .B(n2880), .Y(n1087) );
  INVX1 U2387 ( .A(n2796), .Y(n2778) );
  INVX1 U2388 ( .A(reset), .Y(n2796) );
  INVX1 U2389 ( .A(EN), .Y(n2827) );
  INVX1 U2390 ( .A(WE), .Y(n2844) );
  INVX1 U2391 ( .A(n84), .Y(n2871) );
  INVX1 U2392 ( .A(n2773), .Y(n88) );
  INVX1 U2393 ( .A(n1092), .Y(n2884) );
  INVX1 U2394 ( .A(n85), .Y(n2968) );
  INVX1 U2395 ( .A(n2577), .Y(n2882) );
  INVX1 U2396 ( .A(n2533), .Y(n2883) );
  INVX1 U2397 ( .A(n2774), .Y(n87) );
  INVX1 U2398 ( .A(n2660), .Y(n2983) );
  INVX1 U2399 ( .A(n2661), .Y(n2980) );
  INVX1 U2400 ( .A(n2593), .Y(n2977) );
  INVX1 U2401 ( .A(n2659), .Y(n2974) );
  INVX1 U2402 ( .A(n2658), .Y(n2969) );
  INVX1 U2403 ( .A(n2732), .Y(n2888) );
  INVX1 U2404 ( .A(n2731), .Y(n2876) );
  INVX1 U2405 ( .A(n2543), .Y(n2849) );
  INVX1 U2406 ( .A(n2736), .Y(n2982) );
  INVX1 U2407 ( .A(n2738), .Y(n2979) );
  INVX1 U2408 ( .A(n2737), .Y(n2976) );
  INVX1 U2409 ( .A(n2735), .Y(n2973) );
  INVX1 U2410 ( .A(n2734), .Y(n2970) );
  INVX1 U2411 ( .A(n2664), .Y(n2887) );
  INVX1 U2412 ( .A(n2663), .Y(n2875) );
  INVX1 U2413 ( .A(n2596), .Y(n2845) );
  INVX1 U2414 ( .A(n2617), .Y(n2946) );
  INVX1 U2415 ( .A(n2589), .Y(n2981) );
  INVX1 U2416 ( .A(n2590), .Y(n2978) );
  INVX1 U2417 ( .A(n2657), .Y(n2975) );
  INVX1 U2418 ( .A(n2588), .Y(n2972) );
  INVX1 U2419 ( .A(n2587), .Y(n2971) );
  INVX1 U2420 ( .A(n2542), .Y(n2886) );
  INVX1 U2421 ( .A(n2541), .Y(n2872) );
  INVX1 U2422 ( .A(n2504), .Y(n2850) );
  INVX1 U2423 ( .A(n86), .Y(n2885) );
  INVX1 U2424 ( .A(n2128), .Y(n2848) );
  INVX1 U2425 ( .A(n2080), .Y(n2929) );
  INVX1 U2426 ( .A(n2079), .Y(n2930) );
  INVX1 U2427 ( .A(n2703), .Y(n2938) );
  INVX1 U2428 ( .A(n2618), .Y(n2880) );
  INVX1 U2429 ( .A(n2689), .Y(n2945) );
  INVX1 U2430 ( .A(n2698), .Y(n2941) );
  INVX1 U2431 ( .A(n2687), .Y(n2943) );
  INVX1 U2432 ( .A(n2686), .Y(n2942) );
  INVX1 U2433 ( .A(n2688), .Y(n2944) );
  INVX1 U2434 ( .A(n2694), .Y(n2879) );
  INVX1 U2435 ( .A(n2693), .Y(n2878) );
  INVX1 U2436 ( .A(n2075), .Y(n2937) );
  INVX1 U2437 ( .A(n2076), .Y(n2936) );
  INVX1 U2438 ( .A(n2077), .Y(n2935) );
  INVX1 U2439 ( .A(n2078), .Y(n2934) );
  INVX1 U2440 ( .A(n2081), .Y(n2928) );
  MUX2X1 U2441 ( .B(n2756), .A(n2757), .S(n85), .Y(n2755) );
  MUX2X1 U2442 ( .B(n2759), .A(n2760), .S(n85), .Y(n2758) );
  MUX2X1 U2443 ( .B(n2762), .A(n2763), .S(n85), .Y(n2761) );
  MUX2X1 U2444 ( .B(n2765), .A(n2766), .S(n85), .Y(n2764) );
  MUX2X1 U2445 ( .B(n2768), .A(n2769), .S(n85), .Y(n2767) );
  MUX2X1 U2446 ( .B(n2771), .A(n2772), .S(n85), .Y(n2770) );
  MUX2X1 U2447 ( .B(n2663), .A(n2734), .S(n84), .Y(n2757) );
  MUX2X1 U2448 ( .B(n2735), .A(n2664), .S(n84), .Y(n2756) );
  MUX2X1 U2449 ( .B(n2737), .A(n2738), .S(n84), .Y(n2760) );
  MUX2X1 U2450 ( .B(n2596), .A(n2736), .S(n84), .Y(n2759) );
  MUX2X1 U2451 ( .B(n2758), .A(n2755), .S(n86), .Y(n89) );
  MUX2X1 U2452 ( .B(n2731), .A(n2658), .S(n84), .Y(n2763) );
  MUX2X1 U2453 ( .B(n2659), .A(n2732), .S(n84), .Y(n2762) );
  MUX2X1 U2454 ( .B(n2593), .A(n2661), .S(n84), .Y(n2766) );
  MUX2X1 U2455 ( .B(n2543), .A(n2660), .S(n84), .Y(n2765) );
  MUX2X1 U2456 ( .B(n2764), .A(n2761), .S(n86), .Y(n2773) );
  MUX2X1 U2457 ( .B(n2541), .A(n2587), .S(n84), .Y(n2769) );
  MUX2X1 U2458 ( .B(n2588), .A(n2542), .S(n84), .Y(n2768) );
  MUX2X1 U2459 ( .B(n2657), .A(n2590), .S(n84), .Y(n2772) );
  MUX2X1 U2460 ( .B(n2504), .A(n2589), .S(n84), .Y(n2771) );
  MUX2X1 U2461 ( .B(n2770), .A(n2767), .S(n86), .Y(n2774) );
  MUX2X1 U2462 ( .B(n2984), .A(n2558), .S(n2989), .Y(n252) );
  XOR2X1 U2463 ( .A(n2987), .B(n2988), .Y(n251) );
  XOR2X1 U2464 ( .A(n2823), .B(n236), .Y(n2988) );
  XOR2X1 U2465 ( .A(n235), .B(n233), .Y(n250) );
  XOR2X1 U2466 ( .A(n2818), .B(n2815), .Y(n236) );
  AOI21X1 U2467 ( .A(n2991), .B(DIN[7]), .C(n2992), .Y(n2990) );
  XOR2X1 U2468 ( .A(DIN[7]), .B(n2991), .Y(n235) );
  XOR2X1 U2469 ( .A(DIN[4]), .B(n238), .Y(n2991) );
  AOI21X1 U2470 ( .A(n2994), .B(DIN[3]), .C(n2995), .Y(n2993) );
  XOR2X1 U2471 ( .A(DIN[3]), .B(n2994), .Y(n238) );
  XOR2X1 U2472 ( .A(DIN[6]), .B(DIN[5]), .Y(n2994) );
  AOI21X1 U2473 ( .A(n2997), .B(DIN[0]), .C(n2998), .Y(n2996) );
  XOR2X1 U2474 ( .A(DIN[0]), .B(n2997), .Y(n233) );
  XOR2X1 U2475 ( .A(DIN[1]), .B(DIN[2]), .Y(n2997) );
endmodule


/////////////////////////////////////////////////////////////////
//       testbench: tb.v
/////////////////////////////////////////////////////////////////
`timescale 1ns/10ps
module tb;
integer  a;
integer  b;
initial
begin
a = 3; b = 4;
#5;
a = #5 b + 1;
b <= a + 3;
#10 $stop;
end
endmodule


module lifo ( push, pop, reset, clk, din, empty, full, dout );
  input [15:0] din;
  output [15:0] dout;
  input push, pop, reset, clk;
  output empty, full;
  wire   n34, n35, n36, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727;
  wire   [127:0] mem;

  DFFPOSX1 ptr_reg_0_ ( .D(n383), .CLK(clk), .Q(n34) );
  DFFPOSX1 ptr_reg_1_ ( .D(n408), .CLK(clk), .Q(n35) );
  DFFPOSX1 empty_reg ( .D(n380), .CLK(clk), .Q(empty) );
  DFFPOSX1 dout_reg_0_ ( .D(n687), .CLK(clk), .Q(dout[0]) );
  DFFPOSX1 dout_reg_1_ ( .D(n688), .CLK(clk), .Q(dout[1]) );
  DFFPOSX1 dout_reg_2_ ( .D(n689), .CLK(clk), .Q(dout[2]) );
  DFFPOSX1 dout_reg_3_ ( .D(n690), .CLK(clk), .Q(dout[3]) );
  DFFPOSX1 dout_reg_4_ ( .D(n691), .CLK(clk), .Q(dout[4]) );
  DFFPOSX1 dout_reg_5_ ( .D(n692), .CLK(clk), .Q(dout[5]) );
  DFFPOSX1 dout_reg_6_ ( .D(n693), .CLK(clk), .Q(dout[6]) );
  DFFPOSX1 dout_reg_7_ ( .D(n694), .CLK(clk), .Q(dout[7]) );
  DFFPOSX1 dout_reg_8_ ( .D(n695), .CLK(clk), .Q(dout[8]) );
  DFFPOSX1 dout_reg_9_ ( .D(n696), .CLK(clk), .Q(dout[9]) );
  DFFPOSX1 dout_reg_10_ ( .D(n697), .CLK(clk), .Q(dout[10]) );
  DFFPOSX1 dout_reg_11_ ( .D(n698), .CLK(clk), .Q(dout[11]) );
  DFFPOSX1 dout_reg_12_ ( .D(n699), .CLK(clk), .Q(dout[12]) );
  DFFPOSX1 dout_reg_13_ ( .D(n700), .CLK(clk), .Q(dout[13]) );
  DFFPOSX1 dout_reg_14_ ( .D(n701), .CLK(clk), .Q(dout[14]) );
  DFFPOSX1 dout_reg_15_ ( .D(n702), .CLK(clk), .Q(dout[15]) );
  DFFPOSX1 ptr_reg_2_ ( .D(n382), .CLK(clk), .Q(n36) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n364), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n365), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n366), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n367), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n368), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n369), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n370), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n371), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n372), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n373), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n374), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n375), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n376), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n377), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n378), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n379), .CLK(clk), .Q(mem[0]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n300), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n301), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n302), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n303), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n304), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n305), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n306), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n307), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n308), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n309), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n310), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n311), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n312), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n313), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n314), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n315), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n348), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n349), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n350), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n351), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n352), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n353), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n354), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n355), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n356), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n357), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n358), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n359), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n360), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n361), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n362), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n363), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n332), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n333), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n334), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n335), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n336), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n337), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n338), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n339), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n340), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n341), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n342), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n343), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n344), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n345), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n346), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n347), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n268), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n269), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n270), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n271), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n272), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n273), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n274), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n275), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n276), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n277), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n278), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n279), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n280), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n281), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n282), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n283), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n252), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n253), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n254), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n255), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n256), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n257), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n258), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n259), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n260), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n261), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n262), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n263), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n264), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n265), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n266), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n267), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n316), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n317), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n318), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n319), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n320), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n321), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n322), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n323), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n324), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n325), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n326), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n327), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n328), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n329), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n330), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n331), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n284), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n285), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n286), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n287), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n288), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n289), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n290), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n291), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n292), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n293), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n294), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n295), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n296), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n297), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n298), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n299), .CLK(clk), .Q(mem[80]) );
  OAI21X1 U55 ( .A(n406), .B(n710), .C(n450), .Y(n252) );
  OAI21X1 U57 ( .A(n406), .B(n711), .C(n538), .Y(n253) );
  OAI21X1 U59 ( .A(n406), .B(n712), .C(n551), .Y(n254) );
  OAI21X1 U61 ( .A(n406), .B(n713), .C(n449), .Y(n255) );
  OAI21X1 U63 ( .A(n406), .B(n714), .C(n448), .Y(n256) );
  OAI21X1 U65 ( .A(n406), .B(n715), .C(n468), .Y(n257) );
  OAI21X1 U67 ( .A(n406), .B(n716), .C(n447), .Y(n258) );
  OAI21X1 U69 ( .A(n406), .B(n717), .C(n446), .Y(n259) );
  OAI21X1 U71 ( .A(n406), .B(n718), .C(n497), .Y(n260) );
  OAI21X1 U73 ( .A(n406), .B(n719), .C(n506), .Y(n261) );
  OAI21X1 U75 ( .A(n406), .B(n720), .C(n478), .Y(n262) );
  OAI21X1 U77 ( .A(n406), .B(n721), .C(n488), .Y(n263) );
  OAI21X1 U79 ( .A(n406), .B(n722), .C(n539), .Y(n264) );
  OAI21X1 U81 ( .A(n406), .B(n723), .C(n552), .Y(n265) );
  OAI21X1 U83 ( .A(n406), .B(n724), .C(n515), .Y(n266) );
  OAI21X1 U85 ( .A(n406), .B(n725), .C(n526), .Y(n267) );
  NAND3X1 U87 ( .A(n179), .B(n36), .C(n707), .Y(n55) );
  OAI21X1 U88 ( .A(n710), .B(n684), .C(n536), .Y(n268) );
  OAI21X1 U90 ( .A(n711), .B(n684), .C(n549), .Y(n269) );
  OAI21X1 U92 ( .A(n712), .B(n684), .C(n445), .Y(n270) );
  OAI21X1 U94 ( .A(n713), .B(n684), .C(n444), .Y(n271) );
  OAI21X1 U96 ( .A(n714), .B(n684), .C(n467), .Y(n272) );
  OAI21X1 U98 ( .A(n715), .B(n684), .C(n443), .Y(n273) );
  OAI21X1 U100 ( .A(n716), .B(n684), .C(n442), .Y(n274) );
  OAI21X1 U102 ( .A(n717), .B(n684), .C(n441), .Y(n275) );
  OAI21X1 U104 ( .A(n718), .B(n684), .C(n505), .Y(n276) );
  OAI21X1 U106 ( .A(n719), .B(n684), .C(n496), .Y(n277) );
  OAI21X1 U108 ( .A(n720), .B(n684), .C(n487), .Y(n278) );
  OAI21X1 U110 ( .A(n721), .B(n684), .C(n477), .Y(n279) );
  OAI21X1 U112 ( .A(n722), .B(n684), .C(n550), .Y(n280) );
  OAI21X1 U114 ( .A(n723), .B(n684), .C(n537), .Y(n281) );
  OAI21X1 U116 ( .A(n724), .B(n684), .C(n525), .Y(n282) );
  OAI21X1 U118 ( .A(n725), .B(n684), .C(n514), .Y(n283) );
  OAI21X1 U121 ( .A(n710), .B(n405), .C(n518), .Y(n284) );
  OAI21X1 U123 ( .A(n711), .B(n405), .C(n529), .Y(n285) );
  OAI21X1 U125 ( .A(n712), .B(n405), .C(n440), .Y(n286) );
  OAI21X1 U127 ( .A(n713), .B(n405), .C(n439), .Y(n287) );
  OAI21X1 U129 ( .A(n714), .B(n405), .C(n438), .Y(n288) );
  OAI21X1 U131 ( .A(n715), .B(n405), .C(n437), .Y(n289) );
  OAI21X1 U133 ( .A(n716), .B(n405), .C(n436), .Y(n290) );
  OAI21X1 U135 ( .A(n717), .B(n405), .C(n470), .Y(n291) );
  OAI21X1 U137 ( .A(n718), .B(n405), .C(n480), .Y(n292) );
  OAI21X1 U139 ( .A(n719), .B(n405), .C(n490), .Y(n293) );
  OAI21X1 U141 ( .A(n720), .B(n405), .C(n499), .Y(n294) );
  OAI21X1 U143 ( .A(n721), .B(n405), .C(n508), .Y(n295) );
  OAI21X1 U145 ( .A(n722), .B(n405), .C(n519), .Y(n296) );
  OAI21X1 U147 ( .A(n723), .B(n405), .C(n530), .Y(n297) );
  OAI21X1 U149 ( .A(n724), .B(n405), .C(n541), .Y(n298) );
  OAI21X1 U151 ( .A(n725), .B(n405), .C(n554), .Y(n299) );
  NAND3X1 U153 ( .A(n705), .B(n685), .C(n36), .Y(n105) );
  OAI21X1 U154 ( .A(n123), .B(n710), .C(n435), .Y(n300) );
  OAI21X1 U156 ( .A(n123), .B(n711), .C(n464), .Y(n301) );
  OAI21X1 U158 ( .A(n123), .B(n712), .C(n510), .Y(n302) );
  OAI21X1 U160 ( .A(n123), .B(n713), .C(n521), .Y(n303) );
  OAI21X1 U162 ( .A(n123), .B(n714), .C(n532), .Y(n304) );
  OAI21X1 U164 ( .A(n123), .B(n715), .C(n545), .Y(n305) );
  OAI21X1 U166 ( .A(n123), .B(n716), .C(n434), .Y(n306) );
  OAI21X1 U168 ( .A(n123), .B(n717), .C(n433), .Y(n307) );
  OAI21X1 U170 ( .A(n123), .B(n718), .C(n533), .Y(n308) );
  OAI21X1 U172 ( .A(n123), .B(n719), .C(n546), .Y(n309) );
  OAI21X1 U174 ( .A(n123), .B(n720), .C(n511), .Y(n310) );
  OAI21X1 U176 ( .A(n123), .B(n721), .C(n522), .Y(n311) );
  OAI21X1 U178 ( .A(n123), .B(n722), .C(n493), .Y(n312) );
  OAI21X1 U180 ( .A(n123), .B(n723), .C(n502), .Y(n313) );
  OAI21X1 U182 ( .A(n123), .B(n724), .C(n472), .Y(n314) );
  OAI21X1 U184 ( .A(n123), .B(n725), .C(n482), .Y(n315) );
  NAND3X1 U186 ( .A(n707), .B(n34), .C(n160), .Y(n141) );
  NAND3X1 U187 ( .A(n706), .B(n36), .C(n248), .Y(n140) );
  OAI21X1 U188 ( .A(n710), .B(n683), .C(n527), .Y(n316) );
  OAI21X1 U190 ( .A(n711), .B(n683), .C(n516), .Y(n317) );
  OAI21X1 U192 ( .A(n712), .B(n683), .C(n432), .Y(n318) );
  OAI21X1 U194 ( .A(n713), .B(n683), .C(n431), .Y(n319) );
  OAI21X1 U196 ( .A(n714), .B(n683), .C(n430), .Y(n320) );
  OAI21X1 U198 ( .A(n715), .B(n683), .C(n429), .Y(n321) );
  OAI21X1 U200 ( .A(n716), .B(n683), .C(n469), .Y(n322) );
  OAI21X1 U202 ( .A(n717), .B(n683), .C(n428), .Y(n323) );
  OAI21X1 U204 ( .A(n718), .B(n683), .C(n489), .Y(n324) );
  OAI21X1 U206 ( .A(n719), .B(n683), .C(n479), .Y(n325) );
  OAI21X1 U208 ( .A(n720), .B(n683), .C(n507), .Y(n326) );
  OAI21X1 U210 ( .A(n721), .B(n683), .C(n498), .Y(n327) );
  OAI21X1 U212 ( .A(n722), .B(n683), .C(n528), .Y(n328) );
  OAI21X1 U214 ( .A(n723), .B(n683), .C(n517), .Y(n329) );
  OAI21X1 U216 ( .A(n724), .B(n683), .C(n553), .Y(n330) );
  OAI21X1 U218 ( .A(n725), .B(n683), .C(n540), .Y(n331) );
  AOI22X1 U221 ( .A(n707), .B(n686), .C(n706), .D(n34), .Y(n159) );
  OAI21X1 U222 ( .A(n710), .B(n682), .C(n475), .Y(n332) );
  OAI21X1 U224 ( .A(n711), .B(n682), .C(n485), .Y(n333) );
  OAI21X1 U226 ( .A(n712), .B(n682), .C(n427), .Y(n334) );
  OAI21X1 U228 ( .A(n713), .B(n682), .C(n466), .Y(n335) );
  OAI21X1 U230 ( .A(n714), .B(n682), .C(n426), .Y(n336) );
  OAI21X1 U232 ( .A(n715), .B(n682), .C(n425), .Y(n337) );
  OAI21X1 U234 ( .A(n716), .B(n682), .C(n424), .Y(n338) );
  OAI21X1 U236 ( .A(n717), .B(n682), .C(n423), .Y(n339) );
  OAI21X1 U238 ( .A(n718), .B(n682), .C(n513), .Y(n340) );
  OAI21X1 U240 ( .A(n719), .B(n682), .C(n524), .Y(n341) );
  OAI21X1 U242 ( .A(n720), .B(n682), .C(n535), .Y(n342) );
  OAI21X1 U244 ( .A(n721), .B(n682), .C(n548), .Y(n343) );
  OAI21X1 U246 ( .A(n722), .B(n682), .C(n476), .Y(n344) );
  OAI21X1 U248 ( .A(n723), .B(n682), .C(n486), .Y(n345) );
  OAI21X1 U250 ( .A(n724), .B(n682), .C(n495), .Y(n346) );
  OAI21X1 U252 ( .A(n725), .B(n682), .C(n504), .Y(n347) );
  AOI22X1 U255 ( .A(n180), .B(n707), .C(n706), .D(n179), .Y(n178) );
  OAI21X1 U256 ( .A(n404), .B(n710), .C(n465), .Y(n348) );
  OAI21X1 U258 ( .A(n404), .B(n711), .C(n473), .Y(n349) );
  OAI21X1 U260 ( .A(n404), .B(n712), .C(n483), .Y(n350) );
  OAI21X1 U262 ( .A(n404), .B(n713), .C(n422), .Y(n351) );
  OAI21X1 U264 ( .A(n404), .B(n714), .C(n421), .Y(n352) );
  OAI21X1 U266 ( .A(n404), .B(n715), .C(n420), .Y(n353) );
  OAI21X1 U268 ( .A(n404), .B(n716), .C(n419), .Y(n354) );
  OAI21X1 U270 ( .A(n404), .B(n717), .C(n418), .Y(n355) );
  OAI21X1 U272 ( .A(n404), .B(n718), .C(n523), .Y(n356) );
  OAI21X1 U274 ( .A(n404), .B(n719), .C(n512), .Y(n357) );
  OAI21X1 U276 ( .A(n404), .B(n720), .C(n547), .Y(n358) );
  OAI21X1 U278 ( .A(n404), .B(n721), .C(n534), .Y(n359) );
  OAI21X1 U280 ( .A(n404), .B(n722), .C(n484), .Y(n360) );
  OAI21X1 U282 ( .A(n404), .B(n723), .C(n474), .Y(n361) );
  OAI21X1 U284 ( .A(n404), .B(n724), .C(n503), .Y(n362) );
  OAI21X1 U286 ( .A(n404), .B(n725), .C(n494), .Y(n363) );
  AOI21X1 U288 ( .A(n707), .B(n237), .C(n198), .Y(n181) );
  NOR3X1 U289 ( .A(n557), .B(n36), .C(n543), .Y(n198) );
  NAND3X1 U290 ( .A(n726), .B(n709), .C(n201), .Y(n200) );
  OAI21X1 U291 ( .A(n710), .B(n681), .C(n491), .Y(n364) );
  OAI21X1 U293 ( .A(n711), .B(n681), .C(n500), .Y(n365) );
  OAI21X1 U295 ( .A(n712), .B(n681), .C(n463), .Y(n366) );
  OAI21X1 U297 ( .A(n713), .B(n681), .C(n417), .Y(n367) );
  OAI21X1 U299 ( .A(n714), .B(n681), .C(n416), .Y(n368) );
  OAI21X1 U301 ( .A(n715), .B(n681), .C(n415), .Y(n369) );
  OAI21X1 U303 ( .A(n716), .B(n681), .C(n414), .Y(n370) );
  OAI21X1 U305 ( .A(n717), .B(n681), .C(n413), .Y(n371) );
  OAI21X1 U307 ( .A(n718), .B(n681), .C(n544), .Y(n372) );
  OAI21X1 U309 ( .A(n719), .B(n681), .C(n531), .Y(n373) );
  OAI21X1 U311 ( .A(n720), .B(n681), .C(n520), .Y(n374) );
  OAI21X1 U313 ( .A(n721), .B(n681), .C(n509), .Y(n375) );
  OAI21X1 U315 ( .A(n722), .B(n681), .C(n501), .Y(n376) );
  OAI21X1 U317 ( .A(n723), .B(n681), .C(n492), .Y(n377) );
  OAI21X1 U319 ( .A(n724), .B(n681), .C(n481), .Y(n378) );
  OAI21X1 U321 ( .A(n725), .B(n681), .C(n471), .Y(n379) );
  NAND3X1 U324 ( .A(n201), .B(n709), .C(empty), .Y(n199) );
  AOI22X1 U325 ( .A(dout[15]), .B(n680), .C(n64), .D(n220), .Y(n219) );
  AOI22X1 U326 ( .A(dout[14]), .B(n680), .C(n65), .D(n220), .Y(n221) );
  AOI22X1 U327 ( .A(dout[13]), .B(n680), .C(n66), .D(n220), .Y(n222) );
  AOI22X1 U328 ( .A(dout[12]), .B(n680), .C(n67), .D(n220), .Y(n223) );
  AOI22X1 U329 ( .A(dout[11]), .B(n680), .C(n68), .D(n220), .Y(n224) );
  AOI22X1 U330 ( .A(dout[10]), .B(n680), .C(n69), .D(n220), .Y(n225) );
  AOI22X1 U331 ( .A(dout[9]), .B(n680), .C(n70), .D(n220), .Y(n226) );
  AOI22X1 U332 ( .A(dout[8]), .B(n680), .C(n71), .D(n220), .Y(n227) );
  AOI22X1 U333 ( .A(dout[7]), .B(n679), .C(n72), .D(n220), .Y(n228) );
  AOI22X1 U334 ( .A(dout[6]), .B(n679), .C(n73), .D(n220), .Y(n229) );
  AOI22X1 U335 ( .A(dout[5]), .B(n679), .C(n74), .D(n220), .Y(n230) );
  AOI22X1 U336 ( .A(dout[4]), .B(n679), .C(n75), .D(n220), .Y(n231) );
  AOI22X1 U337 ( .A(dout[3]), .B(n679), .C(n76), .D(n220), .Y(n232) );
  AOI22X1 U338 ( .A(dout[2]), .B(n679), .C(n77), .D(n220), .Y(n233) );
  AOI22X1 U339 ( .A(dout[1]), .B(n679), .C(n78), .D(n220), .Y(n234) );
  AOI22X1 U340 ( .A(dout[0]), .B(n679), .C(n79), .D(n220), .Y(n235) );
  OAI21X1 U341 ( .A(n201), .B(n726), .C(n411), .Y(n380) );
  AOI21X1 U342 ( .A(n703), .B(n237), .C(reset), .Y(n236) );
  NAND3X1 U343 ( .A(n451), .B(n453), .C(n455), .Y(n381) );
  NAND3X1 U345 ( .A(n220), .B(n460), .C(n242), .Y(n239) );
  NAND3X1 U346 ( .A(n461), .B(n458), .C(n462), .Y(n238) );
  OAI21X1 U350 ( .A(n452), .B(n727), .C(n410), .Y(n382) );
  NAND3X1 U351 ( .A(n247), .B(n461), .C(n462), .Y(n246) );
  OAI21X1 U352 ( .A(n686), .B(n556), .C(n727), .Y(n247) );
  AOI21X1 U354 ( .A(n220), .B(n542), .C(n459), .Y(n245) );
  OAI21X1 U356 ( .A(n686), .B(n460), .C(n412), .Y(n383) );
  NAND3X1 U359 ( .A(n461), .B(n709), .C(n454), .Y(n241) );
  NOR3X1 U361 ( .A(full), .B(pop), .C(n708), .Y(n201) );
  NAND3X1 U365 ( .A(n726), .B(n708), .C(pop), .Y(n251) );
  NOR3X1 U366 ( .A(n685), .B(n686), .C(n727), .Y(full) );
  AND2X1 U367 ( .A(n703), .B(n457), .Y(n243) );
  AND2X1 U368 ( .A(n407), .B(n409), .Y(n123) );
  AND2X1 U369 ( .A(n456), .B(n557), .Y(n242) );
  BUFX2 U370 ( .A(n235), .Y(n384) );
  BUFX2 U371 ( .A(n234), .Y(n385) );
  BUFX2 U372 ( .A(n233), .Y(n386) );
  BUFX2 U373 ( .A(n232), .Y(n387) );
  BUFX2 U374 ( .A(n231), .Y(n388) );
  BUFX2 U375 ( .A(n230), .Y(n389) );
  BUFX2 U376 ( .A(n229), .Y(n390) );
  BUFX2 U377 ( .A(n228), .Y(n391) );
  BUFX2 U378 ( .A(n227), .Y(n392) );
  BUFX2 U379 ( .A(n226), .Y(n393) );
  BUFX2 U380 ( .A(n225), .Y(n394) );
  BUFX2 U381 ( .A(n224), .Y(n395) );
  BUFX2 U382 ( .A(n223), .Y(n396) );
  BUFX2 U383 ( .A(n222), .Y(n397) );
  BUFX2 U384 ( .A(n221), .Y(n398) );
  BUFX2 U385 ( .A(n219), .Y(n399) );
  BUFX2 U386 ( .A(n178), .Y(n400) );
  BUFX2 U387 ( .A(n159), .Y(n401) );
  BUFX2 U388 ( .A(n251), .Y(n402) );
  BUFX2 U389 ( .A(n200), .Y(n403) );
  BUFX2 U390 ( .A(n181), .Y(n404) );
  BUFX2 U391 ( .A(n105), .Y(n405) );
  BUFX2 U392 ( .A(n55), .Y(n406) );
  BUFX2 U393 ( .A(n140), .Y(n407) );
  BUFX2 U394 ( .A(n381), .Y(n408) );
  BUFX2 U395 ( .A(n141), .Y(n409) );
  BUFX2 U396 ( .A(n246), .Y(n410) );
  BUFX2 U397 ( .A(n236), .Y(n411) );
  AND2X1 U398 ( .A(n462), .B(n686), .Y(n249) );
  INVX1 U399 ( .A(n249), .Y(n412) );
  AND2X1 U400 ( .A(mem[8]), .B(n681), .Y(n210) );
  INVX1 U401 ( .A(n210), .Y(n413) );
  AND2X1 U402 ( .A(mem[9]), .B(n681), .Y(n209) );
  INVX1 U403 ( .A(n209), .Y(n414) );
  AND2X1 U404 ( .A(mem[10]), .B(n681), .Y(n208) );
  INVX1 U405 ( .A(n208), .Y(n415) );
  AND2X1 U406 ( .A(mem[11]), .B(n681), .Y(n207) );
  INVX1 U407 ( .A(n207), .Y(n416) );
  AND2X1 U408 ( .A(mem[12]), .B(n681), .Y(n206) );
  INVX1 U409 ( .A(n206), .Y(n417) );
  AND2X1 U410 ( .A(mem[24]), .B(n404), .Y(n189) );
  INVX1 U411 ( .A(n189), .Y(n418) );
  AND2X1 U412 ( .A(mem[25]), .B(n404), .Y(n188) );
  INVX1 U413 ( .A(n188), .Y(n419) );
  AND2X1 U414 ( .A(mem[26]), .B(n404), .Y(n187) );
  INVX1 U415 ( .A(n187), .Y(n420) );
  AND2X1 U416 ( .A(mem[27]), .B(n404), .Y(n186) );
  INVX1 U417 ( .A(n186), .Y(n421) );
  AND2X1 U418 ( .A(mem[28]), .B(n404), .Y(n185) );
  INVX1 U419 ( .A(n185), .Y(n422) );
  AND2X1 U420 ( .A(mem[40]), .B(n682), .Y(n169) );
  INVX1 U421 ( .A(n169), .Y(n423) );
  AND2X1 U422 ( .A(mem[41]), .B(n682), .Y(n168) );
  INVX1 U423 ( .A(n168), .Y(n424) );
  AND2X1 U424 ( .A(mem[42]), .B(n682), .Y(n167) );
  INVX1 U425 ( .A(n167), .Y(n425) );
  AND2X1 U426 ( .A(mem[43]), .B(n682), .Y(n166) );
  INVX1 U427 ( .A(n166), .Y(n426) );
  AND2X1 U428 ( .A(mem[45]), .B(n682), .Y(n164) );
  INVX1 U429 ( .A(n164), .Y(n427) );
  AND2X1 U430 ( .A(mem[56]), .B(n683), .Y(n150) );
  INVX1 U431 ( .A(n150), .Y(n428) );
  AND2X1 U432 ( .A(mem[58]), .B(n683), .Y(n148) );
  INVX1 U433 ( .A(n148), .Y(n429) );
  AND2X1 U434 ( .A(mem[59]), .B(n683), .Y(n147) );
  INVX1 U435 ( .A(n147), .Y(n430) );
  AND2X1 U436 ( .A(mem[60]), .B(n683), .Y(n146) );
  INVX1 U437 ( .A(n146), .Y(n431) );
  AND2X1 U438 ( .A(mem[61]), .B(n683), .Y(n145) );
  INVX1 U439 ( .A(n145), .Y(n432) );
  AND2X1 U440 ( .A(mem[72]), .B(n123), .Y(n131) );
  INVX1 U441 ( .A(n131), .Y(n433) );
  AND2X1 U442 ( .A(mem[73]), .B(n123), .Y(n130) );
  INVX1 U443 ( .A(n130), .Y(n434) );
  AND2X1 U444 ( .A(mem[79]), .B(n123), .Y(n124) );
  INVX1 U445 ( .A(n124), .Y(n435) );
  AND2X1 U446 ( .A(mem[89]), .B(n405), .Y(n112) );
  INVX1 U447 ( .A(n112), .Y(n436) );
  AND2X1 U448 ( .A(mem[90]), .B(n405), .Y(n111) );
  INVX1 U449 ( .A(n111), .Y(n437) );
  AND2X1 U450 ( .A(mem[91]), .B(n405), .Y(n110) );
  INVX1 U451 ( .A(n110), .Y(n438) );
  AND2X1 U452 ( .A(mem[92]), .B(n405), .Y(n109) );
  INVX1 U453 ( .A(n109), .Y(n439) );
  AND2X1 U454 ( .A(mem[93]), .B(n405), .Y(n108) );
  INVX1 U455 ( .A(n108), .Y(n440) );
  AND2X1 U456 ( .A(mem[104]), .B(n684), .Y(n96) );
  INVX1 U457 ( .A(n96), .Y(n441) );
  AND2X1 U458 ( .A(mem[105]), .B(n684), .Y(n95) );
  INVX1 U459 ( .A(n95), .Y(n442) );
  AND2X1 U460 ( .A(mem[106]), .B(n684), .Y(n94) );
  INVX1 U461 ( .A(n94), .Y(n443) );
  AND2X1 U462 ( .A(mem[108]), .B(n684), .Y(n92) );
  INVX1 U463 ( .A(n92), .Y(n444) );
  AND2X1 U464 ( .A(mem[109]), .B(n684), .Y(n91) );
  INVX1 U465 ( .A(n91), .Y(n445) );
  AND2X1 U466 ( .A(mem[120]), .B(n406), .Y(n63) );
  INVX1 U467 ( .A(n63), .Y(n446) );
  AND2X1 U468 ( .A(mem[121]), .B(n406), .Y(n62) );
  INVX1 U469 ( .A(n62), .Y(n447) );
  AND2X1 U470 ( .A(mem[123]), .B(n406), .Y(n60) );
  INVX1 U471 ( .A(n60), .Y(n448) );
  AND2X1 U472 ( .A(mem[124]), .B(n406), .Y(n59) );
  INVX1 U473 ( .A(n59), .Y(n449) );
  AND2X1 U474 ( .A(mem[127]), .B(n406), .Y(n56) );
  INVX1 U475 ( .A(n56), .Y(n450) );
  BUFX2 U476 ( .A(n238), .Y(n451) );
  BUFX2 U477 ( .A(n245), .Y(n452) );
  BUFX2 U478 ( .A(n239), .Y(n453) );
  AND2X1 U479 ( .A(n201), .B(n726), .Y(n250) );
  INVX1 U480 ( .A(n250), .Y(n454) );
  AND2X1 U481 ( .A(n459), .B(n678), .Y(n240) );
  INVX1 U482 ( .A(n240), .Y(n455) );
  AND2X1 U483 ( .A(n678), .B(n686), .Y(n179) );
  INVX1 U484 ( .A(n179), .Y(n456) );
  AND2X1 U485 ( .A(n248), .B(n727), .Y(n237) );
  INVX1 U486 ( .A(n237), .Y(n457) );
  INVX1 U487 ( .A(n242), .Y(n458) );
  INVX1 U488 ( .A(n460), .Y(n459) );
  BUFX2 U489 ( .A(n241), .Y(n460) );
  INVX1 U490 ( .A(n243), .Y(n461) );
  OR2X1 U491 ( .A(n459), .B(reset), .Y(n244) );
  INVX1 U492 ( .A(n244), .Y(n462) );
  AND2X1 U493 ( .A(mem[13]), .B(n681), .Y(n205) );
  INVX1 U494 ( .A(n205), .Y(n463) );
  AND2X1 U495 ( .A(mem[78]), .B(n123), .Y(n125) );
  INVX1 U496 ( .A(n125), .Y(n464) );
  AND2X1 U497 ( .A(mem[31]), .B(n404), .Y(n182) );
  INVX1 U498 ( .A(n182), .Y(n465) );
  AND2X1 U499 ( .A(mem[44]), .B(n682), .Y(n165) );
  INVX1 U500 ( .A(n165), .Y(n466) );
  AND2X1 U501 ( .A(mem[107]), .B(n684), .Y(n93) );
  INVX1 U502 ( .A(n93), .Y(n467) );
  AND2X1 U503 ( .A(mem[122]), .B(n406), .Y(n61) );
  INVX1 U504 ( .A(n61), .Y(n468) );
  AND2X1 U505 ( .A(mem[57]), .B(n683), .Y(n149) );
  INVX1 U506 ( .A(n149), .Y(n469) );
  AND2X1 U507 ( .A(mem[88]), .B(n405), .Y(n114) );
  INVX1 U508 ( .A(n114), .Y(n470) );
  AND2X1 U509 ( .A(mem[0]), .B(n681), .Y(n218) );
  INVX1 U510 ( .A(n218), .Y(n471) );
  AND2X1 U511 ( .A(mem[65]), .B(n123), .Y(n138) );
  INVX1 U512 ( .A(n138), .Y(n472) );
  AND2X1 U513 ( .A(mem[30]), .B(n404), .Y(n183) );
  INVX1 U514 ( .A(n183), .Y(n473) );
  AND2X1 U515 ( .A(mem[18]), .B(n404), .Y(n195) );
  INVX1 U516 ( .A(n195), .Y(n474) );
  AND2X1 U517 ( .A(mem[47]), .B(n682), .Y(n162) );
  INVX1 U518 ( .A(n162), .Y(n475) );
  AND2X1 U519 ( .A(mem[35]), .B(n682), .Y(n174) );
  INVX1 U520 ( .A(n174), .Y(n476) );
  AND2X1 U521 ( .A(mem[100]), .B(n684), .Y(n100) );
  INVX1 U522 ( .A(n100), .Y(n477) );
  AND2X1 U523 ( .A(mem[117]), .B(n406), .Y(n82) );
  INVX1 U524 ( .A(n82), .Y(n478) );
  AND2X1 U525 ( .A(mem[54]), .B(n683), .Y(n152) );
  INVX1 U526 ( .A(n152), .Y(n479) );
  AND2X1 U527 ( .A(mem[87]), .B(n405), .Y(n115) );
  INVX1 U528 ( .A(n115), .Y(n480) );
  AND2X1 U529 ( .A(mem[1]), .B(n681), .Y(n217) );
  INVX1 U530 ( .A(n217), .Y(n481) );
  AND2X1 U531 ( .A(mem[64]), .B(n123), .Y(n139) );
  INVX1 U532 ( .A(n139), .Y(n482) );
  AND2X1 U533 ( .A(mem[29]), .B(n404), .Y(n184) );
  INVX1 U534 ( .A(n184), .Y(n483) );
  AND2X1 U535 ( .A(mem[19]), .B(n404), .Y(n194) );
  INVX1 U536 ( .A(n194), .Y(n484) );
  AND2X1 U537 ( .A(mem[46]), .B(n682), .Y(n163) );
  INVX1 U538 ( .A(n163), .Y(n485) );
  AND2X1 U539 ( .A(mem[34]), .B(n682), .Y(n175) );
  INVX1 U540 ( .A(n175), .Y(n486) );
  AND2X1 U541 ( .A(mem[101]), .B(n684), .Y(n99) );
  INVX1 U542 ( .A(n99), .Y(n487) );
  AND2X1 U543 ( .A(mem[116]), .B(n406), .Y(n83) );
  INVX1 U544 ( .A(n83), .Y(n488) );
  AND2X1 U545 ( .A(mem[55]), .B(n683), .Y(n151) );
  INVX1 U546 ( .A(n151), .Y(n489) );
  AND2X1 U547 ( .A(mem[86]), .B(n405), .Y(n116) );
  INVX1 U548 ( .A(n116), .Y(n490) );
  AND2X1 U549 ( .A(mem[15]), .B(n681), .Y(n203) );
  INVX1 U550 ( .A(n203), .Y(n491) );
  AND2X1 U551 ( .A(mem[2]), .B(n681), .Y(n216) );
  INVX1 U552 ( .A(n216), .Y(n492) );
  AND2X1 U553 ( .A(mem[67]), .B(n123), .Y(n136) );
  INVX1 U554 ( .A(n136), .Y(n493) );
  AND2X1 U555 ( .A(mem[16]), .B(n404), .Y(n197) );
  INVX1 U556 ( .A(n197), .Y(n494) );
  AND2X1 U557 ( .A(mem[33]), .B(n682), .Y(n176) );
  INVX1 U558 ( .A(n176), .Y(n495) );
  AND2X1 U559 ( .A(mem[102]), .B(n684), .Y(n98) );
  INVX1 U560 ( .A(n98), .Y(n496) );
  AND2X1 U561 ( .A(mem[119]), .B(n406), .Y(n80) );
  INVX1 U562 ( .A(n80), .Y(n497) );
  AND2X1 U563 ( .A(mem[52]), .B(n683), .Y(n154) );
  INVX1 U564 ( .A(n154), .Y(n498) );
  AND2X1 U565 ( .A(mem[85]), .B(n405), .Y(n117) );
  INVX1 U566 ( .A(n117), .Y(n499) );
  AND2X1 U567 ( .A(mem[14]), .B(n681), .Y(n204) );
  INVX1 U568 ( .A(n204), .Y(n500) );
  AND2X1 U569 ( .A(mem[3]), .B(n681), .Y(n215) );
  INVX1 U570 ( .A(n215), .Y(n501) );
  AND2X1 U571 ( .A(mem[66]), .B(n123), .Y(n137) );
  INVX1 U572 ( .A(n137), .Y(n502) );
  AND2X1 U573 ( .A(mem[17]), .B(n404), .Y(n196) );
  INVX1 U574 ( .A(n196), .Y(n503) );
  AND2X1 U575 ( .A(mem[32]), .B(n682), .Y(n177) );
  INVX1 U576 ( .A(n177), .Y(n504) );
  AND2X1 U577 ( .A(mem[103]), .B(n684), .Y(n97) );
  INVX1 U578 ( .A(n97), .Y(n505) );
  AND2X1 U579 ( .A(mem[118]), .B(n406), .Y(n81) );
  INVX1 U580 ( .A(n81), .Y(n506) );
  AND2X1 U581 ( .A(mem[53]), .B(n683), .Y(n153) );
  INVX1 U582 ( .A(n153), .Y(n507) );
  AND2X1 U583 ( .A(mem[84]), .B(n405), .Y(n118) );
  INVX1 U584 ( .A(n118), .Y(n508) );
  AND2X1 U585 ( .A(mem[4]), .B(n681), .Y(n214) );
  INVX1 U586 ( .A(n214), .Y(n509) );
  AND2X1 U587 ( .A(mem[77]), .B(n123), .Y(n126) );
  INVX1 U588 ( .A(n126), .Y(n510) );
  AND2X1 U589 ( .A(mem[69]), .B(n123), .Y(n134) );
  INVX1 U590 ( .A(n134), .Y(n511) );
  AND2X1 U591 ( .A(mem[22]), .B(n404), .Y(n191) );
  INVX1 U592 ( .A(n191), .Y(n512) );
  AND2X1 U593 ( .A(mem[39]), .B(n682), .Y(n170) );
  INVX1 U594 ( .A(n170), .Y(n513) );
  AND2X1 U595 ( .A(mem[96]), .B(n684), .Y(n104) );
  INVX1 U596 ( .A(n104), .Y(n514) );
  AND2X1 U597 ( .A(mem[113]), .B(n406), .Y(n86) );
  INVX1 U598 ( .A(n86), .Y(n515) );
  AND2X1 U599 ( .A(mem[62]), .B(n683), .Y(n144) );
  INVX1 U600 ( .A(n144), .Y(n516) );
  AND2X1 U601 ( .A(mem[50]), .B(n683), .Y(n156) );
  INVX1 U602 ( .A(n156), .Y(n517) );
  AND2X1 U603 ( .A(mem[95]), .B(n405), .Y(n106) );
  INVX1 U604 ( .A(n106), .Y(n518) );
  AND2X1 U605 ( .A(mem[83]), .B(n405), .Y(n119) );
  INVX1 U606 ( .A(n119), .Y(n519) );
  AND2X1 U607 ( .A(mem[5]), .B(n681), .Y(n213) );
  INVX1 U608 ( .A(n213), .Y(n520) );
  AND2X1 U609 ( .A(mem[76]), .B(n123), .Y(n127) );
  INVX1 U610 ( .A(n127), .Y(n521) );
  AND2X1 U611 ( .A(mem[68]), .B(n123), .Y(n135) );
  INVX1 U612 ( .A(n135), .Y(n522) );
  AND2X1 U613 ( .A(mem[23]), .B(n404), .Y(n190) );
  INVX1 U614 ( .A(n190), .Y(n523) );
  AND2X1 U615 ( .A(mem[38]), .B(n682), .Y(n171) );
  INVX1 U616 ( .A(n171), .Y(n524) );
  AND2X1 U617 ( .A(mem[97]), .B(n684), .Y(n103) );
  INVX1 U618 ( .A(n103), .Y(n525) );
  AND2X1 U619 ( .A(mem[112]), .B(n406), .Y(n87) );
  INVX1 U620 ( .A(n87), .Y(n526) );
  AND2X1 U621 ( .A(mem[63]), .B(n683), .Y(n143) );
  INVX1 U622 ( .A(n143), .Y(n527) );
  AND2X1 U623 ( .A(mem[51]), .B(n683), .Y(n155) );
  INVX1 U624 ( .A(n155), .Y(n528) );
  AND2X1 U625 ( .A(mem[94]), .B(n405), .Y(n107) );
  INVX1 U626 ( .A(n107), .Y(n529) );
  AND2X1 U627 ( .A(mem[82]), .B(n405), .Y(n120) );
  INVX1 U628 ( .A(n120), .Y(n530) );
  AND2X1 U629 ( .A(mem[6]), .B(n681), .Y(n212) );
  INVX1 U630 ( .A(n212), .Y(n531) );
  AND2X1 U631 ( .A(mem[75]), .B(n123), .Y(n128) );
  INVX1 U632 ( .A(n128), .Y(n532) );
  AND2X1 U633 ( .A(mem[71]), .B(n123), .Y(n132) );
  INVX1 U634 ( .A(n132), .Y(n533) );
  AND2X1 U635 ( .A(mem[20]), .B(n404), .Y(n193) );
  INVX1 U636 ( .A(n193), .Y(n534) );
  AND2X1 U637 ( .A(mem[37]), .B(n682), .Y(n172) );
  INVX1 U638 ( .A(n172), .Y(n535) );
  AND2X1 U639 ( .A(mem[111]), .B(n684), .Y(n89) );
  INVX1 U640 ( .A(n89), .Y(n536) );
  AND2X1 U641 ( .A(mem[98]), .B(n684), .Y(n102) );
  INVX1 U642 ( .A(n102), .Y(n537) );
  AND2X1 U643 ( .A(mem[126]), .B(n406), .Y(n57) );
  INVX1 U644 ( .A(n57), .Y(n538) );
  AND2X1 U645 ( .A(mem[115]), .B(n406), .Y(n84) );
  INVX1 U646 ( .A(n84), .Y(n539) );
  AND2X1 U647 ( .A(mem[48]), .B(n683), .Y(n158) );
  INVX1 U648 ( .A(n158), .Y(n540) );
  AND2X1 U649 ( .A(mem[81]), .B(n405), .Y(n121) );
  INVX1 U650 ( .A(n121), .Y(n541) );
  AND2X1 U651 ( .A(n685), .B(n686), .Y(n248) );
  INVX1 U652 ( .A(n248), .Y(n542) );
  BUFX2 U653 ( .A(n199), .Y(n543) );
  AND2X1 U654 ( .A(mem[7]), .B(n681), .Y(n211) );
  INVX1 U655 ( .A(n211), .Y(n544) );
  AND2X1 U656 ( .A(mem[74]), .B(n123), .Y(n129) );
  INVX1 U657 ( .A(n129), .Y(n545) );
  AND2X1 U658 ( .A(mem[70]), .B(n123), .Y(n133) );
  INVX1 U659 ( .A(n133), .Y(n546) );
  AND2X1 U660 ( .A(mem[21]), .B(n404), .Y(n192) );
  INVX1 U661 ( .A(n192), .Y(n547) );
  AND2X1 U662 ( .A(mem[36]), .B(n682), .Y(n173) );
  INVX1 U663 ( .A(n173), .Y(n548) );
  AND2X1 U664 ( .A(mem[110]), .B(n684), .Y(n90) );
  INVX1 U665 ( .A(n90), .Y(n549) );
  AND2X1 U666 ( .A(mem[99]), .B(n684), .Y(n101) );
  INVX1 U667 ( .A(n101), .Y(n550) );
  AND2X1 U668 ( .A(mem[125]), .B(n406), .Y(n58) );
  INVX1 U669 ( .A(n58), .Y(n551) );
  AND2X1 U670 ( .A(mem[114]), .B(n406), .Y(n85) );
  INVX1 U671 ( .A(n85), .Y(n552) );
  AND2X1 U672 ( .A(mem[49]), .B(n683), .Y(n157) );
  INVX1 U673 ( .A(n157), .Y(n553) );
  AND2X1 U674 ( .A(mem[80]), .B(n405), .Y(n122) );
  INVX1 U675 ( .A(n122), .Y(n554) );
  AND2X1 U676 ( .A(n703), .B(n709), .Y(n220) );
  INVX1 U677 ( .A(n220), .Y(n555) );
  AND2X1 U678 ( .A(n678), .B(n727), .Y(n160) );
  INVX1 U679 ( .A(n160), .Y(n556) );
  AND2X1 U680 ( .A(n34), .B(n685), .Y(n180) );
  INVX1 U681 ( .A(n180), .Y(n557) );
  INVX1 U682 ( .A(n558), .Y(n683) );
  INVX1 U683 ( .A(n559), .Y(n681) );
  INVX1 U684 ( .A(n686), .Y(n674) );
  INVX1 U685 ( .A(n686), .Y(n675) );
  INVX1 U686 ( .A(n686), .Y(n676) );
  INVX1 U687 ( .A(n686), .Y(n677) );
  INVX1 U688 ( .A(n685), .Y(n678) );
  BUFX2 U689 ( .A(n555), .Y(n680) );
  AND2X1 U690 ( .A(n160), .B(n705), .Y(n558) );
  AND2X1 U691 ( .A(n237), .B(n706), .Y(n559) );
  BUFX2 U692 ( .A(n555), .Y(n679) );
  INVX1 U693 ( .A(n560), .Y(n682) );
  INVX1 U694 ( .A(n400), .Y(n704) );
  AND2X1 U695 ( .A(n704), .B(n727), .Y(n560) );
  INVX1 U696 ( .A(n543), .Y(n706) );
  INVX1 U697 ( .A(n403), .Y(n707) );
  INVX1 U698 ( .A(n561), .Y(n684) );
  INVX1 U699 ( .A(n401), .Y(n705) );
  INVX1 U700 ( .A(n36), .Y(n727) );
  INVX1 U701 ( .A(din[0]), .Y(n725) );
  INVX1 U702 ( .A(din[1]), .Y(n724) );
  INVX1 U703 ( .A(din[2]), .Y(n723) );
  INVX1 U704 ( .A(din[3]), .Y(n722) );
  INVX1 U705 ( .A(din[4]), .Y(n721) );
  INVX1 U706 ( .A(din[5]), .Y(n720) );
  INVX1 U707 ( .A(din[6]), .Y(n719) );
  INVX1 U708 ( .A(din[7]), .Y(n718) );
  INVX1 U709 ( .A(din[8]), .Y(n717) );
  INVX1 U710 ( .A(din[9]), .Y(n716) );
  INVX1 U711 ( .A(din[10]), .Y(n715) );
  INVX1 U712 ( .A(din[11]), .Y(n714) );
  INVX1 U713 ( .A(din[12]), .Y(n713) );
  INVX1 U714 ( .A(din[13]), .Y(n712) );
  INVX1 U715 ( .A(din[14]), .Y(n711) );
  INVX1 U716 ( .A(din[15]), .Y(n710) );
  AND2X1 U717 ( .A(n36), .B(n704), .Y(n561) );
  INVX1 U718 ( .A(n402), .Y(n703) );
  INVX1 U719 ( .A(n34), .Y(n686) );
  INVX1 U720 ( .A(n399), .Y(n702) );
  INVX1 U721 ( .A(n673), .Y(n64) );
  INVX1 U722 ( .A(n398), .Y(n701) );
  INVX1 U723 ( .A(n672), .Y(n65) );
  INVX1 U724 ( .A(n397), .Y(n700) );
  INVX1 U725 ( .A(n671), .Y(n66) );
  INVX1 U726 ( .A(n396), .Y(n699) );
  INVX1 U727 ( .A(n670), .Y(n67) );
  INVX1 U728 ( .A(n395), .Y(n698) );
  INVX1 U729 ( .A(n669), .Y(n68) );
  INVX1 U730 ( .A(n394), .Y(n697) );
  INVX1 U731 ( .A(n668), .Y(n69) );
  INVX1 U732 ( .A(n393), .Y(n696) );
  INVX1 U733 ( .A(n667), .Y(n70) );
  INVX1 U734 ( .A(n392), .Y(n695) );
  INVX1 U735 ( .A(n666), .Y(n71) );
  INVX1 U736 ( .A(n391), .Y(n694) );
  INVX1 U737 ( .A(n665), .Y(n72) );
  INVX1 U738 ( .A(n390), .Y(n693) );
  INVX1 U739 ( .A(n664), .Y(n73) );
  INVX1 U740 ( .A(n389), .Y(n692) );
  INVX1 U741 ( .A(n663), .Y(n74) );
  INVX1 U742 ( .A(n388), .Y(n691) );
  INVX1 U743 ( .A(n662), .Y(n75) );
  INVX1 U744 ( .A(n387), .Y(n690) );
  INVX1 U745 ( .A(n661), .Y(n76) );
  INVX1 U746 ( .A(n386), .Y(n689) );
  INVX1 U747 ( .A(n660), .Y(n77) );
  INVX1 U748 ( .A(n385), .Y(n688) );
  INVX1 U749 ( .A(n659), .Y(n78) );
  INVX1 U750 ( .A(n384), .Y(n687) );
  INVX1 U751 ( .A(n658), .Y(n79) );
  INVX1 U752 ( .A(n35), .Y(n685) );
  INVX1 U753 ( .A(reset), .Y(n709) );
  INVX1 U754 ( .A(push), .Y(n708) );
  INVX1 U755 ( .A(empty), .Y(n726) );
  MUX2X1 U756 ( .B(n563), .A(n564), .S(n678), .Y(n562) );
  MUX2X1 U757 ( .B(n566), .A(n567), .S(n678), .Y(n565) );
  MUX2X1 U758 ( .B(n569), .A(n570), .S(n678), .Y(n568) );
  MUX2X1 U759 ( .B(n572), .A(n573), .S(n678), .Y(n571) );
  MUX2X1 U760 ( .B(n575), .A(n576), .S(n678), .Y(n574) );
  MUX2X1 U761 ( .B(n578), .A(n579), .S(n678), .Y(n577) );
  MUX2X1 U762 ( .B(n581), .A(n582), .S(n678), .Y(n580) );
  MUX2X1 U763 ( .B(n584), .A(n585), .S(n678), .Y(n583) );
  MUX2X1 U764 ( .B(n587), .A(n588), .S(n678), .Y(n586) );
  MUX2X1 U765 ( .B(n590), .A(n591), .S(n678), .Y(n589) );
  MUX2X1 U766 ( .B(n593), .A(n594), .S(n678), .Y(n592) );
  MUX2X1 U767 ( .B(n596), .A(n597), .S(n678), .Y(n595) );
  MUX2X1 U768 ( .B(n599), .A(n600), .S(n678), .Y(n598) );
  MUX2X1 U769 ( .B(n602), .A(n603), .S(n678), .Y(n601) );
  MUX2X1 U770 ( .B(n605), .A(n606), .S(n678), .Y(n604) );
  MUX2X1 U771 ( .B(n608), .A(n609), .S(n678), .Y(n607) );
  MUX2X1 U772 ( .B(n611), .A(n612), .S(n678), .Y(n610) );
  MUX2X1 U773 ( .B(n614), .A(n615), .S(n678), .Y(n613) );
  MUX2X1 U774 ( .B(n617), .A(n618), .S(n678), .Y(n616) );
  MUX2X1 U775 ( .B(n620), .A(n621), .S(n678), .Y(n619) );
  MUX2X1 U776 ( .B(n623), .A(n624), .S(n678), .Y(n622) );
  MUX2X1 U777 ( .B(n626), .A(n627), .S(n678), .Y(n625) );
  MUX2X1 U778 ( .B(n629), .A(n630), .S(n678), .Y(n628) );
  MUX2X1 U779 ( .B(n632), .A(n633), .S(n678), .Y(n631) );
  MUX2X1 U780 ( .B(n635), .A(n636), .S(n678), .Y(n634) );
  MUX2X1 U781 ( .B(n638), .A(n639), .S(n678), .Y(n637) );
  MUX2X1 U782 ( .B(n641), .A(n642), .S(n678), .Y(n640) );
  MUX2X1 U783 ( .B(n644), .A(n645), .S(n678), .Y(n643) );
  MUX2X1 U784 ( .B(n647), .A(n648), .S(n678), .Y(n646) );
  MUX2X1 U785 ( .B(n650), .A(n651), .S(n678), .Y(n649) );
  MUX2X1 U786 ( .B(n653), .A(n654), .S(n678), .Y(n652) );
  MUX2X1 U787 ( .B(n656), .A(n657), .S(n678), .Y(n655) );
  MUX2X1 U788 ( .B(mem[96]), .A(mem[112]), .S(n677), .Y(n564) );
  MUX2X1 U789 ( .B(mem[64]), .A(mem[80]), .S(n677), .Y(n563) );
  MUX2X1 U790 ( .B(mem[32]), .A(mem[48]), .S(n677), .Y(n567) );
  MUX2X1 U791 ( .B(mem[0]), .A(mem[16]), .S(n677), .Y(n566) );
  MUX2X1 U792 ( .B(n565), .A(n562), .S(n36), .Y(n658) );
  MUX2X1 U793 ( .B(mem[97]), .A(mem[113]), .S(n677), .Y(n570) );
  MUX2X1 U794 ( .B(mem[65]), .A(mem[81]), .S(n677), .Y(n569) );
  MUX2X1 U795 ( .B(mem[33]), .A(mem[49]), .S(n677), .Y(n573) );
  MUX2X1 U796 ( .B(mem[1]), .A(mem[17]), .S(n677), .Y(n572) );
  MUX2X1 U797 ( .B(n571), .A(n568), .S(n36), .Y(n659) );
  MUX2X1 U798 ( .B(mem[98]), .A(mem[114]), .S(n677), .Y(n576) );
  MUX2X1 U799 ( .B(mem[66]), .A(mem[82]), .S(n677), .Y(n575) );
  MUX2X1 U800 ( .B(mem[34]), .A(mem[50]), .S(n677), .Y(n579) );
  MUX2X1 U801 ( .B(mem[2]), .A(mem[18]), .S(n677), .Y(n578) );
  MUX2X1 U802 ( .B(n577), .A(n574), .S(n36), .Y(n660) );
  MUX2X1 U803 ( .B(mem[99]), .A(mem[115]), .S(n676), .Y(n582) );
  MUX2X1 U804 ( .B(mem[67]), .A(mem[83]), .S(n676), .Y(n581) );
  MUX2X1 U805 ( .B(mem[35]), .A(mem[51]), .S(n676), .Y(n585) );
  MUX2X1 U806 ( .B(mem[3]), .A(mem[19]), .S(n676), .Y(n584) );
  MUX2X1 U807 ( .B(n583), .A(n580), .S(n36), .Y(n661) );
  MUX2X1 U808 ( .B(mem[100]), .A(mem[116]), .S(n676), .Y(n588) );
  MUX2X1 U809 ( .B(mem[68]), .A(mem[84]), .S(n676), .Y(n587) );
  MUX2X1 U810 ( .B(mem[36]), .A(mem[52]), .S(n676), .Y(n591) );
  MUX2X1 U811 ( .B(mem[4]), .A(mem[20]), .S(n676), .Y(n590) );
  MUX2X1 U812 ( .B(n589), .A(n586), .S(n36), .Y(n662) );
  MUX2X1 U813 ( .B(mem[101]), .A(mem[117]), .S(n676), .Y(n594) );
  MUX2X1 U814 ( .B(mem[69]), .A(mem[85]), .S(n676), .Y(n593) );
  MUX2X1 U815 ( .B(mem[37]), .A(mem[53]), .S(n676), .Y(n597) );
  MUX2X1 U816 ( .B(mem[5]), .A(mem[21]), .S(n676), .Y(n596) );
  MUX2X1 U817 ( .B(n595), .A(n592), .S(n36), .Y(n663) );
  MUX2X1 U818 ( .B(mem[102]), .A(mem[118]), .S(n675), .Y(n600) );
  MUX2X1 U819 ( .B(mem[70]), .A(mem[86]), .S(n675), .Y(n599) );
  MUX2X1 U820 ( .B(mem[38]), .A(mem[54]), .S(n675), .Y(n603) );
  MUX2X1 U821 ( .B(mem[6]), .A(mem[22]), .S(n675), .Y(n602) );
  MUX2X1 U822 ( .B(n601), .A(n598), .S(n36), .Y(n664) );
  MUX2X1 U823 ( .B(mem[103]), .A(mem[119]), .S(n675), .Y(n606) );
  MUX2X1 U824 ( .B(mem[71]), .A(mem[87]), .S(n675), .Y(n605) );
  MUX2X1 U825 ( .B(mem[39]), .A(mem[55]), .S(n675), .Y(n609) );
  MUX2X1 U826 ( .B(mem[7]), .A(mem[23]), .S(n675), .Y(n608) );
  MUX2X1 U827 ( .B(n607), .A(n604), .S(n36), .Y(n665) );
  MUX2X1 U828 ( .B(mem[104]), .A(mem[120]), .S(n675), .Y(n612) );
  MUX2X1 U829 ( .B(mem[72]), .A(mem[88]), .S(n675), .Y(n611) );
  MUX2X1 U830 ( .B(mem[40]), .A(mem[56]), .S(n675), .Y(n615) );
  MUX2X1 U831 ( .B(mem[8]), .A(mem[24]), .S(n675), .Y(n614) );
  MUX2X1 U832 ( .B(n613), .A(n610), .S(n36), .Y(n666) );
  MUX2X1 U833 ( .B(mem[105]), .A(mem[121]), .S(n674), .Y(n618) );
  MUX2X1 U834 ( .B(mem[73]), .A(mem[89]), .S(n674), .Y(n617) );
  MUX2X1 U835 ( .B(mem[41]), .A(mem[57]), .S(n674), .Y(n621) );
  MUX2X1 U836 ( .B(mem[9]), .A(mem[25]), .S(n674), .Y(n620) );
  MUX2X1 U837 ( .B(n619), .A(n616), .S(n36), .Y(n667) );
  MUX2X1 U838 ( .B(mem[106]), .A(mem[122]), .S(n674), .Y(n624) );
  MUX2X1 U839 ( .B(mem[74]), .A(mem[90]), .S(n674), .Y(n623) );
  MUX2X1 U840 ( .B(mem[42]), .A(mem[58]), .S(n674), .Y(n627) );
  MUX2X1 U841 ( .B(mem[10]), .A(mem[26]), .S(n674), .Y(n626) );
  MUX2X1 U842 ( .B(n625), .A(n622), .S(n36), .Y(n668) );
  MUX2X1 U843 ( .B(mem[107]), .A(mem[123]), .S(n674), .Y(n630) );
  MUX2X1 U844 ( .B(mem[75]), .A(mem[91]), .S(n674), .Y(n629) );
  MUX2X1 U845 ( .B(mem[43]), .A(mem[59]), .S(n674), .Y(n633) );
  MUX2X1 U846 ( .B(mem[11]), .A(mem[27]), .S(n674), .Y(n632) );
  MUX2X1 U847 ( .B(n631), .A(n628), .S(n36), .Y(n669) );
  MUX2X1 U848 ( .B(mem[108]), .A(mem[124]), .S(n674), .Y(n636) );
  MUX2X1 U849 ( .B(mem[76]), .A(mem[92]), .S(n677), .Y(n635) );
  MUX2X1 U850 ( .B(mem[44]), .A(mem[60]), .S(n676), .Y(n639) );
  MUX2X1 U851 ( .B(mem[12]), .A(mem[28]), .S(n675), .Y(n638) );
  MUX2X1 U852 ( .B(n637), .A(n634), .S(n36), .Y(n670) );
  MUX2X1 U853 ( .B(mem[109]), .A(mem[125]), .S(n677), .Y(n642) );
  MUX2X1 U854 ( .B(mem[77]), .A(mem[93]), .S(n676), .Y(n641) );
  MUX2X1 U855 ( .B(mem[45]), .A(mem[61]), .S(n675), .Y(n645) );
  MUX2X1 U856 ( .B(mem[13]), .A(mem[29]), .S(n674), .Y(n644) );
  MUX2X1 U857 ( .B(n643), .A(n640), .S(n36), .Y(n671) );
  MUX2X1 U858 ( .B(mem[110]), .A(mem[126]), .S(n676), .Y(n648) );
  MUX2X1 U859 ( .B(mem[78]), .A(mem[94]), .S(n675), .Y(n647) );
  MUX2X1 U860 ( .B(mem[46]), .A(mem[62]), .S(n674), .Y(n651) );
  MUX2X1 U861 ( .B(mem[14]), .A(mem[30]), .S(n677), .Y(n650) );
  MUX2X1 U862 ( .B(n649), .A(n646), .S(n36), .Y(n672) );
  MUX2X1 U863 ( .B(mem[111]), .A(mem[127]), .S(n676), .Y(n654) );
  MUX2X1 U864 ( .B(mem[79]), .A(mem[95]), .S(n677), .Y(n653) );
  MUX2X1 U865 ( .B(mem[47]), .A(mem[63]), .S(n674), .Y(n657) );
  MUX2X1 U866 ( .B(mem[15]), .A(mem[31]), .S(n675), .Y(n656) );
  MUX2X1 U867 ( .B(n655), .A(n652), .S(n36), .Y(n673) );
endmodule



module FIFO_DEPTH_P25_WIDTH16 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, net263, net264,
         net265;
  wire   [4:0] wr_ptr;
  wire   [4:0] rd_ptr;
  wire   [511:0] mem;
  tri   clk;
  tri   reset;
  tri   get;
  tri   [15:0] data_out;
  assign full = fillcount[5];

  \**SEQGEN**  mem_reg_31__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[511]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[510]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[509]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[508]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[507]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[506]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[505]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[504]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[503]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[502]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[501]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[500]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[499]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[498]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[497]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[496]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_30__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[495]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[494]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[493]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[492]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[491]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[490]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[489]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[488]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[487]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[486]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[485]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[484]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[483]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[482]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[481]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[480]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_29__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[479]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[478]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[477]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[476]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[475]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[474]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[473]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[472]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[471]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[470]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[469]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[468]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[467]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[466]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[465]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[464]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_28__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[463]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[462]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[461]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[460]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[459]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[458]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[457]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[456]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[455]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[454]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[453]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[452]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[451]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[450]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[449]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[448]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_27__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[447]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[446]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[445]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[444]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[443]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[442]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[441]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[440]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[439]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[438]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[437]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[436]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[435]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[434]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[433]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[432]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_26__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[431]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[430]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[429]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[428]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[427]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[426]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[425]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[424]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[423]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[422]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[421]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[420]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[419]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[418]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[417]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[416]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_25__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[415]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[414]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[413]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[412]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[411]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[410]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[409]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[408]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[407]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[406]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[405]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[404]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[403]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[402]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[401]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[400]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_24__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[399]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[398]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[397]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[396]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[395]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[394]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[393]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[392]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[391]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[390]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[389]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[388]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[387]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[386]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[385]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[384]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_23__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[383]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[382]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[381]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[380]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[379]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[378]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[377]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[376]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[375]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[374]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[373]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[372]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[371]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[370]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[369]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[368]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_22__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[367]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[366]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[365]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[364]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[363]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[362]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[361]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[360]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[359]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[358]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[357]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[356]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[355]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[354]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[353]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[352]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_21__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[351]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[350]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[349]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[348]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[347]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[346]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[345]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[344]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[343]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[342]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[341]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[340]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[339]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[338]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[337]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[336]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_20__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[335]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[334]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[333]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[332]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[331]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[330]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[329]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[328]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[327]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[326]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[325]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[324]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[323]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[322]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[321]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[320]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_19__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[319]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[318]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[317]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[316]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[315]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[314]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[313]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[312]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[311]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[310]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[309]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[308]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[307]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[306]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[305]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[304]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_18__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[303]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[302]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[301]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[300]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[299]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[298]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[297]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[296]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[295]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[294]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[293]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[292]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[291]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[290]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[289]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[288]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_17__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[287]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[286]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[285]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[284]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[283]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[282]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[281]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[280]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[279]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[278]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[277]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[276]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[275]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[274]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[273]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[272]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_16__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[271]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[270]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[269]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[268]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[267]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[266]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[265]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[264]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[263]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[262]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[261]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[260]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[259]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[258]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[257]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[256]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_15__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_14__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_13__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_12__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_11__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_10__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_9__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_8__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_7__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_6__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[99]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[98]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[97]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[96]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N90) );
  \**SEQGEN**  mem_reg_5__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[95]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[94]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[93]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[92]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[91]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[90]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[89]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[88]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[87]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[86]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[85]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[84]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[83]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[82]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[81]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[80]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N89) );
  \**SEQGEN**  mem_reg_4__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[79]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[78]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[77]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[76]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[75]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[74]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[73]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[72]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[71]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[70]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[69]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[68]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[67]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[66]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[65]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[64]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N88) );
  \**SEQGEN**  mem_reg_3__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[63]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[62]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[61]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[60]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[59]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[58]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[57]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[56]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[55]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[54]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[53]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[52]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[51]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[50]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[49]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[48]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N87) );
  \**SEQGEN**  mem_reg_2__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[47]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[46]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[45]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[44]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[43]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[42]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[41]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[40]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[39]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[38]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[37]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[36]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[35]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[34]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[33]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[32]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_1__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_0__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  fillcount_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N83), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N82), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N81), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N80), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N79), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N78), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  rd_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  wr_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  GTECH_OR2 C3419 ( .A(fillcount[4]), .B(fillcount[5]), .Z(N124) );
  GTECH_OR2 C3420 ( .A(fillcount[3]), .B(N124), .Z(N125) );
  GTECH_OR2 C3421 ( .A(fillcount[2]), .B(N125), .Z(N126) );
  GTECH_OR2 C3422 ( .A(fillcount[1]), .B(N126), .Z(N127) );
  GTECH_OR2 C3423 ( .A(fillcount[0]), .B(N127), .Z(N128) );
  GTECH_NOT I_0 ( .A(N128), .Z(empty) );
  ADD_UNS_OP add_33 ( .A(rd_ptr), .B(1'b1), .Z({N40, N39, N38, N37, N36}) );
  ADD_UNS_OP add_32 ( .A(wr_ptr), .B(1'b1), .Z({N35, N34, N33, N32, N31}) );
  GTECH_OR3 C3425 ( .A(reset), .B(N117), .C(N120), .Z(N65) );
  GTECH_OR3 C3440 ( .A(reset), .B(N117), .C(N123), .Z(N71) );
  GTECH_OR3 C3455 ( .A(reset), .B(N120), .C(N123), .Z(N77) );
  ADD_UNS_OP add_37 ( .A(fillcount), .B(1'b1), .Z({N52, N51, N50, N49, N48, 
        N47}) );
  ADD_UNS_OP add_36 ( .A(wr_ptr), .B(1'b1), .Z({N46, N45, N44, N43, N42}) );
  SUB_UNS_OP sub_40 ( .A(fillcount), .B(1'b1), .Z({N64, N63, N62, N61, N60, 
        N59}) );
  ADD_UNS_OP add_39 ( .A(rd_ptr), .B(1'b1), .Z({N58, N57, N56, N55, N54}) );
  GTECH_OR3 C3473 ( .A(reset), .B(N123), .C(N29), .Z(N130) );
  GTECH_AND2 C4497 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N131) );
  GTECH_AND2 C4498 ( .A(N0), .B(wr_ptr[4]), .Z(N132) );
  GTECH_NOT I_1 ( .A(wr_ptr[3]), .Z(N0) );
  GTECH_AND2 C4499 ( .A(wr_ptr[3]), .B(N1), .Z(N133) );
  GTECH_NOT I_2 ( .A(wr_ptr[4]), .Z(N1) );
  GTECH_AND2 C4500 ( .A(N2), .B(N3), .Z(N134) );
  GTECH_NOT I_3 ( .A(wr_ptr[3]), .Z(N2) );
  GTECH_NOT I_4 ( .A(wr_ptr[4]), .Z(N3) );
  GTECH_NOT I_5 ( .A(wr_ptr[2]), .Z(N135) );
  GTECH_AND2 C4502 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N136) );
  GTECH_AND2 C4503 ( .A(N4), .B(wr_ptr[1]), .Z(N137) );
  GTECH_NOT I_6 ( .A(wr_ptr[0]), .Z(N4) );
  GTECH_AND2 C4504 ( .A(wr_ptr[0]), .B(N5), .Z(N138) );
  GTECH_NOT I_7 ( .A(wr_ptr[1]), .Z(N5) );
  GTECH_AND2 C4505 ( .A(N6), .B(N7), .Z(N139) );
  GTECH_NOT I_8 ( .A(wr_ptr[0]), .Z(N6) );
  GTECH_NOT I_9 ( .A(wr_ptr[1]), .Z(N7) );
  GTECH_AND2 C4506 ( .A(wr_ptr[2]), .B(N136), .Z(N140) );
  GTECH_AND2 C4507 ( .A(wr_ptr[2]), .B(N137), .Z(N141) );
  GTECH_AND2 C4508 ( .A(wr_ptr[2]), .B(N138), .Z(N142) );
  GTECH_AND2 C4509 ( .A(wr_ptr[2]), .B(N139), .Z(N143) );
  GTECH_AND2 C4510 ( .A(N135), .B(N136), .Z(N144) );
  GTECH_AND2 C4511 ( .A(N135), .B(N137), .Z(N145) );
  GTECH_AND2 C4512 ( .A(N135), .B(N138), .Z(N146) );
  GTECH_AND2 C4513 ( .A(N135), .B(N139), .Z(N147) );
  GTECH_AND2 C4514 ( .A(N131), .B(N140), .Z(N148) );
  GTECH_AND2 C4515 ( .A(N131), .B(N141), .Z(N149) );
  GTECH_AND2 C4516 ( .A(N131), .B(N142), .Z(N150) );
  GTECH_AND2 C4517 ( .A(N131), .B(N143), .Z(N151) );
  GTECH_AND2 C4518 ( .A(N131), .B(N144), .Z(N152) );
  GTECH_AND2 C4519 ( .A(N131), .B(N145), .Z(N153) );
  GTECH_AND2 C4520 ( .A(N131), .B(N146), .Z(N154) );
  GTECH_AND2 C4521 ( .A(N131), .B(N147), .Z(N155) );
  GTECH_AND2 C4522 ( .A(N132), .B(N140), .Z(N156) );
  GTECH_AND2 C4523 ( .A(N132), .B(N141), .Z(N157) );
  GTECH_AND2 C4524 ( .A(N132), .B(N142), .Z(N158) );
  GTECH_AND2 C4525 ( .A(N132), .B(N143), .Z(N159) );
  GTECH_AND2 C4526 ( .A(N132), .B(N144), .Z(N160) );
  GTECH_AND2 C4527 ( .A(N132), .B(N145), .Z(N161) );
  GTECH_AND2 C4528 ( .A(N132), .B(N146), .Z(N162) );
  GTECH_AND2 C4529 ( .A(N132), .B(N147), .Z(N163) );
  GTECH_AND2 C4530 ( .A(N133), .B(N140), .Z(N164) );
  GTECH_AND2 C4531 ( .A(N133), .B(N141), .Z(N165) );
  GTECH_AND2 C4532 ( .A(N133), .B(N142), .Z(N166) );
  GTECH_AND2 C4533 ( .A(N133), .B(N143), .Z(N167) );
  GTECH_AND2 C4534 ( .A(N133), .B(N144), .Z(N168) );
  GTECH_AND2 C4535 ( .A(N133), .B(N145), .Z(N169) );
  GTECH_AND2 C4536 ( .A(N133), .B(N146), .Z(N170) );
  GTECH_AND2 C4537 ( .A(N133), .B(N147), .Z(N171) );
  GTECH_AND2 C4538 ( .A(N134), .B(N140), .Z(N172) );
  GTECH_AND2 C4539 ( .A(N134), .B(N141), .Z(N173) );
  GTECH_AND2 C4540 ( .A(N134), .B(N142), .Z(N174) );
  GTECH_AND2 C4541 ( .A(N134), .B(N143), .Z(N175) );
  GTECH_AND2 C4542 ( .A(N134), .B(N144), .Z(N176) );
  GTECH_AND2 C4543 ( .A(N134), .B(N145), .Z(N177) );
  GTECH_AND2 C4544 ( .A(N134), .B(N146), .Z(N178) );
  GTECH_AND2 C4545 ( .A(N134), .B(N147), .Z(N179) );
  GTECH_AND2 C4546 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N180) );
  GTECH_AND2 C4547 ( .A(N8), .B(wr_ptr[4]), .Z(N181) );
  GTECH_NOT I_10 ( .A(wr_ptr[3]), .Z(N8) );
  GTECH_AND2 C4548 ( .A(wr_ptr[3]), .B(N9), .Z(N182) );
  GTECH_NOT I_11 ( .A(wr_ptr[4]), .Z(N9) );
  GTECH_AND2 C4549 ( .A(N10), .B(N11), .Z(N183) );
  GTECH_NOT I_12 ( .A(wr_ptr[3]), .Z(N10) );
  GTECH_NOT I_13 ( .A(wr_ptr[4]), .Z(N11) );
  GTECH_AND2 C4551 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N184) );
  GTECH_AND2 C4552 ( .A(N12), .B(wr_ptr[1]), .Z(N185) );
  GTECH_NOT I_14 ( .A(wr_ptr[0]), .Z(N12) );
  GTECH_AND2 C4553 ( .A(wr_ptr[0]), .B(N13), .Z(N186) );
  GTECH_NOT I_15 ( .A(wr_ptr[1]), .Z(N13) );
  GTECH_AND2 C4554 ( .A(N14), .B(N15), .Z(N187) );
  GTECH_NOT I_16 ( .A(wr_ptr[0]), .Z(N14) );
  GTECH_NOT I_17 ( .A(wr_ptr[1]), .Z(N15) );
  GTECH_AND2 C4555 ( .A(wr_ptr[2]), .B(N184), .Z(N188) );
  GTECH_AND2 C4556 ( .A(wr_ptr[2]), .B(N185), .Z(N189) );
  GTECH_AND2 C4557 ( .A(wr_ptr[2]), .B(N186), .Z(N190) );
  GTECH_AND2 C4558 ( .A(wr_ptr[2]), .B(N187), .Z(N191) );
  GTECH_AND2 C4559 ( .A(N135), .B(N184), .Z(N192) );
  GTECH_AND2 C4560 ( .A(N135), .B(N185), .Z(N193) );
  GTECH_AND2 C4561 ( .A(N135), .B(N186), .Z(N194) );
  GTECH_AND2 C4562 ( .A(N135), .B(N187), .Z(N195) );
  GTECH_AND2 C4563 ( .A(N180), .B(N188), .Z(N196) );
  GTECH_AND2 C4564 ( .A(N180), .B(N189), .Z(N197) );
  GTECH_AND2 C4565 ( .A(N180), .B(N190), .Z(N198) );
  GTECH_AND2 C4566 ( .A(N180), .B(N191), .Z(N199) );
  GTECH_AND2 C4567 ( .A(N180), .B(N192), .Z(N200) );
  GTECH_AND2 C4568 ( .A(N180), .B(N193), .Z(N201) );
  GTECH_AND2 C4569 ( .A(N180), .B(N194), .Z(N202) );
  GTECH_AND2 C4570 ( .A(N180), .B(N195), .Z(N203) );
  GTECH_AND2 C4571 ( .A(N181), .B(N188), .Z(N204) );
  GTECH_AND2 C4572 ( .A(N181), .B(N189), .Z(N205) );
  GTECH_AND2 C4573 ( .A(N181), .B(N190), .Z(N206) );
  GTECH_AND2 C4574 ( .A(N181), .B(N191), .Z(N207) );
  GTECH_AND2 C4575 ( .A(N181), .B(N192), .Z(N208) );
  GTECH_AND2 C4576 ( .A(N181), .B(N193), .Z(N209) );
  GTECH_AND2 C4577 ( .A(N181), .B(N194), .Z(N210) );
  GTECH_AND2 C4578 ( .A(N181), .B(N195), .Z(N211) );
  GTECH_AND2 C4579 ( .A(N182), .B(N188), .Z(N212) );
  GTECH_AND2 C4580 ( .A(N182), .B(N189), .Z(N213) );
  GTECH_AND2 C4581 ( .A(N182), .B(N190), .Z(N214) );
  GTECH_AND2 C4582 ( .A(N182), .B(N191), .Z(N215) );
  GTECH_AND2 C4583 ( .A(N182), .B(N192), .Z(N216) );
  GTECH_AND2 C4584 ( .A(N182), .B(N193), .Z(N217) );
  GTECH_AND2 C4585 ( .A(N182), .B(N194), .Z(N218) );
  GTECH_AND2 C4586 ( .A(N182), .B(N195), .Z(N219) );
  GTECH_AND2 C4587 ( .A(N183), .B(N188), .Z(N220) );
  GTECH_AND2 C4588 ( .A(N183), .B(N189), .Z(N221) );
  GTECH_AND2 C4589 ( .A(N183), .B(N190), .Z(N222) );
  GTECH_AND2 C4590 ( .A(N183), .B(N191), .Z(N223) );
  GTECH_AND2 C4591 ( .A(N183), .B(N192), .Z(N224) );
  GTECH_AND2 C4592 ( .A(N183), .B(N193), .Z(N225) );
  GTECH_AND2 C4593 ( .A(N183), .B(N194), .Z(N226) );
  GTECH_AND2 C4594 ( .A(N183), .B(N195), .Z(N227) );
  SELECT_OP C4595 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N35, N34, 
        N33, N32, N31}), .DATA3({N46, N45, N44, N43, N42}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N120), .Z({N70, N69, N68, N67, N66}) );
  GTECH_BUF B_0 ( .A(reset), .Z(N16) );
  SELECT_OP C4596 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N40, N39, 
        N38, N37, N36}), .DATA3({N58, N57, N56, N55, N54}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N123), .Z({N76, N75, N74, N73, N72}) );
  SELECT_OP C4597 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N52, 
        N51, N50, N49, N48, N47}), .DATA3({N64, N63, N62, N61, N60, N59}), 
        .CONTROL1(N16), .CONTROL2(N120), .CONTROL3(N123), .Z({N83, N82, N81, 
        N80, N79, N78}) );
  SELECT_OP C4598 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
        N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
        N171, N172, N173, N174, N175, N176, N177, N178, N179}), .DATA3({N196, 
        N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
        N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
        N221, N222, N223, N224, N225, N226, N227}), .CONTROL1(N17), .CONTROL2(
        N117), .CONTROL3(N120), .Z({N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84}) );
  GTECH_BUF B_1 ( .A(N130), .Z(N17) );
  MUX_OP C4599 ( .D0({mem[0], mem[1], mem[2], mem[3], mem[4], mem[5], mem[6], 
        mem[7], mem[8], mem[9], mem[10], mem[11], mem[12], mem[13], mem[14], 
        mem[15]}), .D1({mem[16], mem[17], mem[18], mem[19], mem[20], mem[21], 
        mem[22], mem[23], mem[24], mem[25], mem[26], mem[27], mem[28], mem[29], 
        mem[30], mem[31]}), .D2({mem[32], mem[33], mem[34], mem[35], mem[36], 
        mem[37], mem[38], mem[39], mem[40], mem[41], mem[42], mem[43], mem[44], 
        mem[45], mem[46], mem[47]}), .D3({mem[48], mem[49], mem[50], mem[51], 
        mem[52], mem[53], mem[54], mem[55], mem[56], mem[57], mem[58], mem[59], 
        mem[60], mem[61], mem[62], mem[63]}), .D4({mem[64], mem[65], mem[66], 
        mem[67], mem[68], mem[69], mem[70], mem[71], mem[72], mem[73], mem[74], 
        mem[75], mem[76], mem[77], mem[78], mem[79]}), .D5({mem[80], mem[81], 
        mem[82], mem[83], mem[84], mem[85], mem[86], mem[87], mem[88], mem[89], 
        mem[90], mem[91], mem[92], mem[93], mem[94], mem[95]}), .D6({mem[96], 
        mem[97], mem[98], mem[99], mem[100], mem[101], mem[102], mem[103], 
        mem[104], mem[105], mem[106], mem[107], mem[108], mem[109], mem[110], 
        mem[111]}), .D7({mem[112], mem[113], mem[114], mem[115], mem[116], 
        mem[117], mem[118], mem[119], mem[120], mem[121], mem[122], mem[123], 
        mem[124], mem[125], mem[126], mem[127]}), .D8({mem[128], mem[129], 
        mem[130], mem[131], mem[132], mem[133], mem[134], mem[135], mem[136], 
        mem[137], mem[138], mem[139], mem[140], mem[141], mem[142], mem[143]}), 
        .D9({mem[144], mem[145], mem[146], mem[147], mem[148], mem[149], 
        mem[150], mem[151], mem[152], mem[153], mem[154], mem[155], mem[156], 
        mem[157], mem[158], mem[159]}), .D10({mem[160], mem[161], mem[162], 
        mem[163], mem[164], mem[165], mem[166], mem[167], mem[168], mem[169], 
        mem[170], mem[171], mem[172], mem[173], mem[174], mem[175]}), .D11({
        mem[176], mem[177], mem[178], mem[179], mem[180], mem[181], mem[182], 
        mem[183], mem[184], mem[185], mem[186], mem[187], mem[188], mem[189], 
        mem[190], mem[191]}), .D12({mem[192], mem[193], mem[194], mem[195], 
        mem[196], mem[197], mem[198], mem[199], mem[200], mem[201], mem[202], 
        mem[203], mem[204], mem[205], mem[206], mem[207]}), .D13({mem[208], 
        mem[209], mem[210], mem[211], mem[212], mem[213], mem[214], mem[215], 
        mem[216], mem[217], mem[218], mem[219], mem[220], mem[221], mem[222], 
        mem[223]}), .D14({mem[224], mem[225], mem[226], mem[227], mem[228], 
        mem[229], mem[230], mem[231], mem[232], mem[233], mem[234], mem[235], 
        mem[236], mem[237], mem[238], mem[239]}), .D15({mem[240], mem[241], 
        mem[242], mem[243], mem[244], mem[245], mem[246], mem[247], mem[248], 
        mem[249], mem[250], mem[251], mem[252], mem[253], mem[254], mem[255]}), 
        .D16({mem[256], mem[257], mem[258], mem[259], mem[260], mem[261], 
        mem[262], mem[263], mem[264], mem[265], mem[266], mem[267], mem[268], 
        mem[269], mem[270], mem[271]}), .D17({mem[272], mem[273], mem[274], 
        mem[275], mem[276], mem[277], mem[278], mem[279], mem[280], mem[281], 
        mem[282], mem[283], mem[284], mem[285], mem[286], mem[287]}), .D18({
        mem[288], mem[289], mem[290], mem[291], mem[292], mem[293], mem[294], 
        mem[295], mem[296], mem[297], mem[298], mem[299], mem[300], mem[301], 
        mem[302], mem[303]}), .D19({mem[304], mem[305], mem[306], mem[307], 
        mem[308], mem[309], mem[310], mem[311], mem[312], mem[313], mem[314], 
        mem[315], mem[316], mem[317], mem[318], mem[319]}), .D20({mem[320], 
        mem[321], mem[322], mem[323], mem[324], mem[325], mem[326], mem[327], 
        mem[328], mem[329], mem[330], mem[331], mem[332], mem[333], mem[334], 
        mem[335]}), .D21({mem[336], mem[337], mem[338], mem[339], mem[340], 
        mem[341], mem[342], mem[343], mem[344], mem[345], mem[346], mem[347], 
        mem[348], mem[349], mem[350], mem[351]}), .D22({mem[352], mem[353], 
        mem[354], mem[355], mem[356], mem[357], mem[358], mem[359], mem[360], 
        mem[361], mem[362], mem[363], mem[364], mem[365], mem[366], mem[367]}), 
        .D23({mem[368], mem[369], mem[370], mem[371], mem[372], mem[373], 
        mem[374], mem[375], mem[376], mem[377], mem[378], mem[379], mem[380], 
        mem[381], mem[382], mem[383]}), .D24({mem[384], mem[385], mem[386], 
        mem[387], mem[388], mem[389], mem[390], mem[391], mem[392], mem[393], 
        mem[394], mem[395], mem[396], mem[397], mem[398], mem[399]}), .D25({
        mem[400], mem[401], mem[402], mem[403], mem[404], mem[405], mem[406], 
        mem[407], mem[408], mem[409], mem[410], mem[411], mem[412], mem[413], 
        mem[414], mem[415]}), .D26({mem[416], mem[417], mem[418], mem[419], 
        mem[420], mem[421], mem[422], mem[423], mem[424], mem[425], mem[426], 
        mem[427], mem[428], mem[429], mem[430], mem[431]}), .D27({mem[432], 
        mem[433], mem[434], mem[435], mem[436], mem[437], mem[438], mem[439], 
        mem[440], mem[441], mem[442], mem[443], mem[444], mem[445], mem[446], 
        mem[447]}), .D28({mem[448], mem[449], mem[450], mem[451], mem[452], 
        mem[453], mem[454], mem[455], mem[456], mem[457], mem[458], mem[459], 
        mem[460], mem[461], mem[462], mem[463]}), .D29({mem[464], mem[465], 
        mem[466], mem[467], mem[468], mem[469], mem[470], mem[471], mem[472], 
        mem[473], mem[474], mem[475], mem[476], mem[477], mem[478], mem[479]}), 
        .D30({mem[480], mem[481], mem[482], mem[483], mem[484], mem[485], 
        mem[486], mem[487], mem[488], mem[489], mem[490], mem[491], mem[492], 
        mem[493], mem[494], mem[495]}), .D31({mem[496], mem[497], mem[498], 
        mem[499], mem[500], mem[501], mem[502], mem[503], mem[504], mem[505], 
        mem[506], mem[507], mem[508], mem[509], mem[510], mem[511]}), .S0(N18), 
        .S1(N19), .S2(N20), .S3(N21), .S4(N22), .Z({data_out[0], data_out[1], 
        data_out[2], data_out[3], data_out[4], data_out[5], data_out[6], 
        data_out[7], data_out[8], data_out[9], data_out[10], data_out[11], 
        data_out[12], data_out[13], data_out[14], data_out[15]}) );
  GTECH_BUF B_2 ( .A(rd_ptr[0]), .Z(N18) );
  GTECH_BUF B_3 ( .A(rd_ptr[1]), .Z(N19) );
  GTECH_BUF B_4 ( .A(rd_ptr[2]), .Z(N20) );
  GTECH_BUF B_5 ( .A(rd_ptr[3]), .Z(N21) );
  GTECH_BUF B_6 ( .A(rd_ptr[4]), .Z(N22) );
  GTECH_AND2 C4602 ( .A(N228), .B(put), .Z(N23) );
  GTECH_NOT I_18 ( .A(fillcount[5]), .Z(N228) );
  GTECH_AND2 C4605 ( .A(N229), .B(get), .Z(N24) );
  GTECH_AND2 C4606 ( .A(N23), .B(N128), .Z(N229) );
  GTECH_AND2 C4607 ( .A(N128), .B(get), .Z(N25) );
  GTECH_OR2 C4612 ( .A(N24), .B(reset), .Z(N26) );
  GTECH_OR2 C4613 ( .A(N23), .B(N26), .Z(N27) );
  GTECH_OR2 C4614 ( .A(N25), .B(N27), .Z(N28) );
  GTECH_NOT I_19 ( .A(N28), .Z(N29) );
  GTECH_BUF B_7 ( .A(N117), .Z(N30) );
  GTECH_BUF B_8 ( .A(N120), .Z(N41) );
  GTECH_BUF B_9 ( .A(N123), .Z(N53) );
  GTECH_NOT I_20 ( .A(reset), .Z(N116) );
  GTECH_AND2 C4684 ( .A(N24), .B(N116), .Z(N117) );
  GTECH_AND2 C4685 ( .A(N30), .B(N116), .Z(net263) );
  GTECH_NOT I_21 ( .A(N24), .Z(N118) );
  GTECH_AND2 C4687 ( .A(N116), .B(N118), .Z(N119) );
  GTECH_AND2 C4688 ( .A(N23), .B(N119), .Z(N120) );
  GTECH_AND2 C4689 ( .A(N41), .B(N119), .Z(net264) );
  GTECH_NOT I_22 ( .A(N23), .Z(N121) );
  GTECH_AND2 C4691 ( .A(N119), .B(N121), .Z(N122) );
  GTECH_AND2 C4692 ( .A(N25), .B(N122), .Z(N123) );
  GTECH_AND2 C4693 ( .A(N53), .B(N122), .Z(net265) );
endmodule


module FIFO_DEPTH_P25_WIDTH34 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [33:0] data_in;
  output [33:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, net342, net343,
         net344;
  wire   [4:0] wr_ptr;
  wire   [4:0] rd_ptr;
  wire   [1087:0] mem;
  tri   clk;
  tri   reset;
  tri   get;
  tri   [33:0] data_out;
  tri   empty;
  assign full = fillcount[5];

  \**SEQGEN**  mem_reg_31__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1087]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1086]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1085]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1084]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1083]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1082]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1081]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1080]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1079]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1078]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1077]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1076]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1075]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1074]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1073]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1072]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1071]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1070]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1069]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1068]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1067]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1066]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1065]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1064]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1063]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1062]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1061]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1060]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1059]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1058]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1057]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1056]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1055]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1054]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_30__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1053]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1052]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1051]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1050]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1049]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1048]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1047]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1046]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1045]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1044]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1043]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1042]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1041]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1040]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1039]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1038]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1037]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1036]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1035]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1034]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1033]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1032]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1031]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1030]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1029]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1028]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1027]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1026]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1025]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1024]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1023]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1022]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1021]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1020]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_29__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1019]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1018]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1017]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1016]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1015]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1014]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1013]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1012]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1011]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1010]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1009]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1008]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1007]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1006]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1005]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1004]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1003]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1002]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1001]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1000]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[999]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[998]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[997]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[996]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[995]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[994]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[993]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[992]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[991]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[990]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[989]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[988]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[987]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[986]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_28__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[985]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[984]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[983]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[982]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[981]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[980]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[979]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[978]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[977]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[976]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[975]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[974]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[973]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[972]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[971]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[970]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[969]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[968]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[967]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[966]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[965]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[964]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[963]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[962]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[961]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[960]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[959]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[958]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[957]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[956]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[955]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[954]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[953]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[952]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_27__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[951]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[950]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[949]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[948]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[947]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[946]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[945]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[944]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[943]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[942]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[941]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[940]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[939]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[938]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[937]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[936]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[935]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[934]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[933]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[932]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[931]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[930]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[929]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[928]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[927]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[926]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[925]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[924]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[923]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[922]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[921]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[920]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[919]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[918]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_26__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[917]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[916]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[915]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[914]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[913]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[912]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[911]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[910]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[909]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[908]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[907]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[906]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[905]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[904]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[903]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[902]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[901]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[900]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[899]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[898]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[897]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[896]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[895]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[894]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[893]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[892]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[891]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[890]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[889]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[888]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[887]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[886]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[885]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[884]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_25__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[883]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[882]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[881]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[880]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[879]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[878]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[877]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[876]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[875]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[874]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[873]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[872]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[871]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[870]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[869]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[868]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[867]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[866]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[865]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[864]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[863]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[862]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[861]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[860]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[859]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[858]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[857]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[856]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[855]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[854]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[853]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[852]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[851]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[850]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_24__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[849]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[848]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[847]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[846]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[845]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[844]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[843]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[842]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[841]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[840]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[839]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[838]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[837]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[836]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[835]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[834]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[833]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[832]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[831]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[830]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[829]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[828]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[827]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[826]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[825]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[824]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[823]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[822]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[821]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[820]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[819]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[818]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[817]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[816]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_23__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[815]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[814]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[813]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[812]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[811]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[810]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[809]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[808]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[807]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[806]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[805]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[804]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[803]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[802]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[801]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[800]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[799]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[798]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[797]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[796]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[795]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[794]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[793]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[792]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[791]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[790]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[789]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[788]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[787]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[786]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[785]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[784]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[783]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[782]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_22__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[781]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[780]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[779]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[778]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[777]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[776]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[775]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[774]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[773]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[772]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[771]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[770]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[769]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[768]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[767]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[766]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[765]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[764]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[763]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[762]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[761]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[760]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[759]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[758]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[757]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[756]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[755]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[754]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[753]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[752]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[751]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[750]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[749]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[748]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_21__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[747]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[746]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[745]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[744]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[743]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[742]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[741]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[740]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[739]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[738]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[737]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[736]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[735]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[734]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[733]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[732]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[731]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[730]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[729]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[728]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[727]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[726]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[725]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[724]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[723]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[722]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[721]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[720]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[719]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[718]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[717]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[716]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[715]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[714]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_20__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[713]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[712]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[711]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[710]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[709]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[708]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[707]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[706]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[705]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[704]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[703]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[702]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[701]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[700]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[699]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[698]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[697]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[696]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[695]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[694]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[693]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[692]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[691]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[690]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[689]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[688]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[687]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[686]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[685]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[684]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[683]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[682]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[681]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[680]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_19__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[679]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[678]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[677]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[676]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[675]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[674]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[673]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[672]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[671]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[670]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[669]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[668]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[667]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[666]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[665]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[664]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[663]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[662]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[661]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[660]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[659]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[658]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[657]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[656]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[655]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[654]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[653]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[652]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[651]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[650]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[649]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[648]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[647]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[646]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_18__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[645]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[644]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[643]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[642]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[641]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[640]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[639]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[638]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[637]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[636]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[635]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[634]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[633]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[632]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[631]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[630]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[629]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[628]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[627]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[626]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[625]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[624]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[623]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[622]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[621]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[620]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[619]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[618]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[617]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[616]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[615]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[614]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[613]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[612]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_17__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[611]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[610]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[609]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[608]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[607]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[606]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[605]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[604]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[603]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[602]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[601]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[600]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[599]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[598]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[597]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[596]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[595]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[594]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[593]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[592]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[591]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[590]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[589]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[588]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[587]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[586]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[585]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[584]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[583]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[582]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[581]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[580]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[579]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[578]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_16__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[577]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[576]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[575]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[574]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[573]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[572]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[571]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[570]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[569]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[568]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[567]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[566]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[565]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[564]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[563]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[562]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[561]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[560]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[559]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[558]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[557]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[556]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[555]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[554]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[553]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[552]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[551]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[550]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[549]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[548]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[547]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[546]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[545]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[544]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_15__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[543]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[542]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[541]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[540]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[539]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[538]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[537]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[536]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[535]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[534]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[533]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[532]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[531]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[530]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[529]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[528]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[527]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[526]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[525]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[524]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[523]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[522]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[521]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[520]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[519]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[518]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[517]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[516]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[515]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[514]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[513]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[512]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[511]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[510]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_14__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[509]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[508]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[507]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[506]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[505]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[504]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[503]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[502]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[501]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[500]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[499]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[498]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[497]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[496]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[495]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[494]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[493]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[492]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[491]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[490]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[489]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[488]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[487]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[486]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[485]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[484]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[483]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[482]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[481]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[480]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[479]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[478]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[477]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[476]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_13__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[475]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[474]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[473]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[472]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[471]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[470]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[469]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[468]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[467]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[466]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[465]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[464]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[463]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[462]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[461]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[460]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[459]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[458]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[457]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[456]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[455]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[454]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[453]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[452]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[451]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[450]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[449]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[448]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[447]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[446]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[445]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[444]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[443]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[442]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_12__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[441]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[440]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[439]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[438]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[437]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[436]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[435]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[434]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[433]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[432]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[431]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[430]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[429]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[428]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[427]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[426]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[425]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[424]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[423]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[422]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[421]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[420]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[419]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[418]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[417]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[416]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[415]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[414]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[413]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[412]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[411]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[410]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[409]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[408]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_11__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[407]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[406]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[405]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[404]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[403]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[402]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[401]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[400]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[399]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[398]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[397]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[396]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[395]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[394]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[393]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[392]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[391]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[390]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[389]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[388]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[387]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[386]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[385]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[384]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[383]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[382]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[381]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[380]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[379]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[378]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[377]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[376]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[375]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[374]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_10__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[373]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[372]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[371]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[370]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[369]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[368]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[367]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[366]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[365]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[364]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[363]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[362]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[361]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[360]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[359]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[358]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[357]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[356]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[355]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[354]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[353]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[352]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[351]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[350]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[349]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[348]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[347]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[346]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[345]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[344]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[343]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[342]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[341]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[340]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_9__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[339]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[338]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[337]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[336]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[335]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[334]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[333]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[332]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[331]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[330]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[329]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[328]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[327]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[326]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[325]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[324]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[323]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[322]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[321]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[320]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[319]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[318]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[317]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[316]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[315]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[314]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[313]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[312]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[311]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[310]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[309]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[308]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[307]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[306]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_8__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[305]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[304]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[303]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[302]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[301]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[300]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[299]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[298]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[297]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[296]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[295]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[294]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[293]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[292]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[291]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[290]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[289]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[288]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[287]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[286]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[285]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[284]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[283]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[282]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[281]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[280]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[279]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[278]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[277]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[276]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[275]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[274]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[273]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[272]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_7__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[271]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[270]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[269]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[268]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[267]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[266]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[265]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[264]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[263]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[262]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[261]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[260]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[259]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[258]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[257]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[256]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_6__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_5__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_4__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_3__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_2__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[99]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[98]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[97]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[96]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[95]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[94]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[93]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[92]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[91]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[90]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[89]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[88]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[87]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[86]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[85]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[84]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[83]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[82]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[81]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[80]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[79]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[78]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[77]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[76]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[75]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[74]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[73]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[72]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[71]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[70]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[69]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[68]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_1__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[67]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[66]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[65]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[64]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[63]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[62]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[61]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[60]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[59]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[58]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[57]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[56]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[55]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[54]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[53]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[52]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[51]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[50]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[49]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[48]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[47]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[46]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[45]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[44]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[43]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[42]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[41]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[40]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[39]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[38]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[37]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[36]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[35]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[34]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_0__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[33]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[32]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  fillcount_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N83), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N82), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N81), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N80), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N79), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N78), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  rd_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  wr_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  GTECH_OR2 C6875 ( .A(fillcount[4]), .B(fillcount[5]), .Z(N124) );
  GTECH_OR2 C6876 ( .A(fillcount[3]), .B(N124), .Z(N125) );
  GTECH_OR2 C6877 ( .A(fillcount[2]), .B(N125), .Z(N126) );
  GTECH_OR2 C6878 ( .A(fillcount[1]), .B(N126), .Z(N127) );
  GTECH_OR2 C6879 ( .A(fillcount[0]), .B(N127), .Z(N128) );
  GTECH_NOT I_0 ( .A(N128), .Z(empty) );
  ADD_UNS_OP add_33 ( .A(rd_ptr), .B(1'b1), .Z({N40, N39, N38, N37, N36}) );
  ADD_UNS_OP add_32 ( .A(wr_ptr), .B(1'b1), .Z({N35, N34, N33, N32, N31}) );
  GTECH_OR3 C6881 ( .A(reset), .B(N117), .C(N120), .Z(N65) );
  GTECH_OR3 C6896 ( .A(reset), .B(N117), .C(N123), .Z(N71) );
  GTECH_OR3 C6911 ( .A(reset), .B(N120), .C(N123), .Z(N77) );
  ADD_UNS_OP add_37 ( .A(fillcount), .B(1'b1), .Z({N52, N51, N50, N49, N48, 
        N47}) );
  ADD_UNS_OP add_36 ( .A(wr_ptr), .B(1'b1), .Z({N46, N45, N44, N43, N42}) );
  SUB_UNS_OP sub_40 ( .A(fillcount), .B(1'b1), .Z({N64, N63, N62, N61, N60, 
        N59}) );
  ADD_UNS_OP add_39 ( .A(rd_ptr), .B(1'b1), .Z({N58, N57, N56, N55, N54}) );
  GTECH_OR3 C6929 ( .A(reset), .B(N123), .C(N29), .Z(N130) );
  GTECH_AND2 C9105 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N131) );
  GTECH_AND2 C9106 ( .A(N0), .B(wr_ptr[4]), .Z(N132) );
  GTECH_NOT I_1 ( .A(wr_ptr[3]), .Z(N0) );
  GTECH_AND2 C9107 ( .A(wr_ptr[3]), .B(N1), .Z(N133) );
  GTECH_NOT I_2 ( .A(wr_ptr[4]), .Z(N1) );
  GTECH_AND2 C9108 ( .A(N2), .B(N3), .Z(N134) );
  GTECH_NOT I_3 ( .A(wr_ptr[3]), .Z(N2) );
  GTECH_NOT I_4 ( .A(wr_ptr[4]), .Z(N3) );
  GTECH_NOT I_5 ( .A(wr_ptr[2]), .Z(N135) );
  GTECH_AND2 C9110 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N136) );
  GTECH_AND2 C9111 ( .A(N4), .B(wr_ptr[1]), .Z(N137) );
  GTECH_NOT I_6 ( .A(wr_ptr[0]), .Z(N4) );
  GTECH_AND2 C9112 ( .A(wr_ptr[0]), .B(N5), .Z(N138) );
  GTECH_NOT I_7 ( .A(wr_ptr[1]), .Z(N5) );
  GTECH_AND2 C9113 ( .A(N6), .B(N7), .Z(N139) );
  GTECH_NOT I_8 ( .A(wr_ptr[0]), .Z(N6) );
  GTECH_NOT I_9 ( .A(wr_ptr[1]), .Z(N7) );
  GTECH_AND2 C9114 ( .A(wr_ptr[2]), .B(N136), .Z(N140) );
  GTECH_AND2 C9115 ( .A(wr_ptr[2]), .B(N137), .Z(N141) );
  GTECH_AND2 C9116 ( .A(wr_ptr[2]), .B(N138), .Z(N142) );
  GTECH_AND2 C9117 ( .A(wr_ptr[2]), .B(N139), .Z(N143) );
  GTECH_AND2 C9118 ( .A(N135), .B(N136), .Z(N144) );
  GTECH_AND2 C9119 ( .A(N135), .B(N137), .Z(N145) );
  GTECH_AND2 C9120 ( .A(N135), .B(N138), .Z(N146) );
  GTECH_AND2 C9121 ( .A(N135), .B(N139), .Z(N147) );
  GTECH_AND2 C9122 ( .A(N131), .B(N140), .Z(N148) );
  GTECH_AND2 C9123 ( .A(N131), .B(N141), .Z(N149) );
  GTECH_AND2 C9124 ( .A(N131), .B(N142), .Z(N150) );
  GTECH_AND2 C9125 ( .A(N131), .B(N143), .Z(N151) );
  GTECH_AND2 C9126 ( .A(N131), .B(N144), .Z(N152) );
  GTECH_AND2 C9127 ( .A(N131), .B(N145), .Z(N153) );
  GTECH_AND2 C9128 ( .A(N131), .B(N146), .Z(N154) );
  GTECH_AND2 C9129 ( .A(N131), .B(N147), .Z(N155) );
  GTECH_AND2 C9130 ( .A(N132), .B(N140), .Z(N156) );
  GTECH_AND2 C9131 ( .A(N132), .B(N141), .Z(N157) );
  GTECH_AND2 C9132 ( .A(N132), .B(N142), .Z(N158) );
  GTECH_AND2 C9133 ( .A(N132), .B(N143), .Z(N159) );
  GTECH_AND2 C9134 ( .A(N132), .B(N144), .Z(N160) );
  GTECH_AND2 C9135 ( .A(N132), .B(N145), .Z(N161) );
  GTECH_AND2 C9136 ( .A(N132), .B(N146), .Z(N162) );
  GTECH_AND2 C9137 ( .A(N132), .B(N147), .Z(N163) );
  GTECH_AND2 C9138 ( .A(N133), .B(N140), .Z(N164) );
  GTECH_AND2 C9139 ( .A(N133), .B(N141), .Z(N165) );
  GTECH_AND2 C9140 ( .A(N133), .B(N142), .Z(N166) );
  GTECH_AND2 C9141 ( .A(N133), .B(N143), .Z(N167) );
  GTECH_AND2 C9142 ( .A(N133), .B(N144), .Z(N168) );
  GTECH_AND2 C9143 ( .A(N133), .B(N145), .Z(N169) );
  GTECH_AND2 C9144 ( .A(N133), .B(N146), .Z(N170) );
  GTECH_AND2 C9145 ( .A(N133), .B(N147), .Z(N171) );
  GTECH_AND2 C9146 ( .A(N134), .B(N140), .Z(N172) );
  GTECH_AND2 C9147 ( .A(N134), .B(N141), .Z(N173) );
  GTECH_AND2 C9148 ( .A(N134), .B(N142), .Z(N174) );
  GTECH_AND2 C9149 ( .A(N134), .B(N143), .Z(N175) );
  GTECH_AND2 C9150 ( .A(N134), .B(N144), .Z(N176) );
  GTECH_AND2 C9151 ( .A(N134), .B(N145), .Z(N177) );
  GTECH_AND2 C9152 ( .A(N134), .B(N146), .Z(N178) );
  GTECH_AND2 C9153 ( .A(N134), .B(N147), .Z(N179) );
  GTECH_AND2 C9154 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N180) );
  GTECH_AND2 C9155 ( .A(N8), .B(wr_ptr[4]), .Z(N181) );
  GTECH_NOT I_10 ( .A(wr_ptr[3]), .Z(N8) );
  GTECH_AND2 C9156 ( .A(wr_ptr[3]), .B(N9), .Z(N182) );
  GTECH_NOT I_11 ( .A(wr_ptr[4]), .Z(N9) );
  GTECH_AND2 C9157 ( .A(N10), .B(N11), .Z(N183) );
  GTECH_NOT I_12 ( .A(wr_ptr[3]), .Z(N10) );
  GTECH_NOT I_13 ( .A(wr_ptr[4]), .Z(N11) );
  GTECH_AND2 C9159 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N184) );
  GTECH_AND2 C9160 ( .A(N12), .B(wr_ptr[1]), .Z(N185) );
  GTECH_NOT I_14 ( .A(wr_ptr[0]), .Z(N12) );
  GTECH_AND2 C9161 ( .A(wr_ptr[0]), .B(N13), .Z(N186) );
  GTECH_NOT I_15 ( .A(wr_ptr[1]), .Z(N13) );
  GTECH_AND2 C9162 ( .A(N14), .B(N15), .Z(N187) );
  GTECH_NOT I_16 ( .A(wr_ptr[0]), .Z(N14) );
  GTECH_NOT I_17 ( .A(wr_ptr[1]), .Z(N15) );
  GTECH_AND2 C9163 ( .A(wr_ptr[2]), .B(N184), .Z(N188) );
  GTECH_AND2 C9164 ( .A(wr_ptr[2]), .B(N185), .Z(N189) );
  GTECH_AND2 C9165 ( .A(wr_ptr[2]), .B(N186), .Z(N190) );
  GTECH_AND2 C9166 ( .A(wr_ptr[2]), .B(N187), .Z(N191) );
  GTECH_AND2 C9167 ( .A(N135), .B(N184), .Z(N192) );
  GTECH_AND2 C9168 ( .A(N135), .B(N185), .Z(N193) );
  GTECH_AND2 C9169 ( .A(N135), .B(N186), .Z(N194) );
  GTECH_AND2 C9170 ( .A(N135), .B(N187), .Z(N195) );
  GTECH_AND2 C9171 ( .A(N180), .B(N188), .Z(N196) );
  GTECH_AND2 C9172 ( .A(N180), .B(N189), .Z(N197) );
  GTECH_AND2 C9173 ( .A(N180), .B(N190), .Z(N198) );
  GTECH_AND2 C9174 ( .A(N180), .B(N191), .Z(N199) );
  GTECH_AND2 C9175 ( .A(N180), .B(N192), .Z(N200) );
  GTECH_AND2 C9176 ( .A(N180), .B(N193), .Z(N201) );
  GTECH_AND2 C9177 ( .A(N180), .B(N194), .Z(N202) );
  GTECH_AND2 C9178 ( .A(N180), .B(N195), .Z(N203) );
  GTECH_AND2 C9179 ( .A(N181), .B(N188), .Z(N204) );
  GTECH_AND2 C9180 ( .A(N181), .B(N189), .Z(N205) );
  GTECH_AND2 C9181 ( .A(N181), .B(N190), .Z(N206) );
  GTECH_AND2 C9182 ( .A(N181), .B(N191), .Z(N207) );
  GTECH_AND2 C9183 ( .A(N181), .B(N192), .Z(N208) );
  GTECH_AND2 C9184 ( .A(N181), .B(N193), .Z(N209) );
  GTECH_AND2 C9185 ( .A(N181), .B(N194), .Z(N210) );
  GTECH_AND2 C9186 ( .A(N181), .B(N195), .Z(N211) );
  GTECH_AND2 C9187 ( .A(N182), .B(N188), .Z(N212) );
  GTECH_AND2 C9188 ( .A(N182), .B(N189), .Z(N213) );
  GTECH_AND2 C9189 ( .A(N182), .B(N190), .Z(N214) );
  GTECH_AND2 C9190 ( .A(N182), .B(N191), .Z(N215) );
  GTECH_AND2 C9191 ( .A(N182), .B(N192), .Z(N216) );
  GTECH_AND2 C9192 ( .A(N182), .B(N193), .Z(N217) );
  GTECH_AND2 C9193 ( .A(N182), .B(N194), .Z(N218) );
  GTECH_AND2 C9194 ( .A(N182), .B(N195), .Z(N219) );
  GTECH_AND2 C9195 ( .A(N183), .B(N188), .Z(N220) );
  GTECH_AND2 C9196 ( .A(N183), .B(N189), .Z(N221) );
  GTECH_AND2 C9197 ( .A(N183), .B(N190), .Z(N222) );
  GTECH_AND2 C9198 ( .A(N183), .B(N191), .Z(N223) );
  GTECH_AND2 C9199 ( .A(N183), .B(N192), .Z(N224) );
  GTECH_AND2 C9200 ( .A(N183), .B(N193), .Z(N225) );
  GTECH_AND2 C9201 ( .A(N183), .B(N194), .Z(N226) );
  GTECH_AND2 C9202 ( .A(N183), .B(N195), .Z(N227) );
  SELECT_OP C9203 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N35, N34, 
        N33, N32, N31}), .DATA3({N46, N45, N44, N43, N42}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N120), .Z({N70, N69, N68, N67, N66}) );
  GTECH_BUF B_0 ( .A(reset), .Z(N16) );
  SELECT_OP C9204 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N40, N39, 
        N38, N37, N36}), .DATA3({N58, N57, N56, N55, N54}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N123), .Z({N76, N75, N74, N73, N72}) );
  SELECT_OP C9205 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N52, 
        N51, N50, N49, N48, N47}), .DATA3({N64, N63, N62, N61, N60, N59}), 
        .CONTROL1(N16), .CONTROL2(N120), .CONTROL3(N123), .Z({N83, N82, N81, 
        N80, N79, N78}) );
  SELECT_OP C9206 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
        N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
        N171, N172, N173, N174, N175, N176, N177, N178, N179}), .DATA3({N196, 
        N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
        N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
        N221, N222, N223, N224, N225, N226, N227}), .CONTROL1(N17), .CONTROL2(
        N117), .CONTROL3(N120), .Z({N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84}) );
  GTECH_BUF B_1 ( .A(N130), .Z(N17) );
  MUX_OP C9207 ( .D0({mem[0], mem[1], mem[2], mem[3], mem[4], mem[5], mem[6], 
        mem[7], mem[8], mem[9], mem[10], mem[11], mem[12], mem[13], mem[14], 
        mem[15], mem[16], mem[17], mem[18], mem[19], mem[20], mem[21], mem[22], 
        mem[23], mem[24], mem[25], mem[26], mem[27], mem[28], mem[29], mem[30], 
        mem[31], mem[32], mem[33]}), .D1({mem[34], mem[35], mem[36], mem[37], 
        mem[38], mem[39], mem[40], mem[41], mem[42], mem[43], mem[44], mem[45], 
        mem[46], mem[47], mem[48], mem[49], mem[50], mem[51], mem[52], mem[53], 
        mem[54], mem[55], mem[56], mem[57], mem[58], mem[59], mem[60], mem[61], 
        mem[62], mem[63], mem[64], mem[65], mem[66], mem[67]}), .D2({mem[68], 
        mem[69], mem[70], mem[71], mem[72], mem[73], mem[74], mem[75], mem[76], 
        mem[77], mem[78], mem[79], mem[80], mem[81], mem[82], mem[83], mem[84], 
        mem[85], mem[86], mem[87], mem[88], mem[89], mem[90], mem[91], mem[92], 
        mem[93], mem[94], mem[95], mem[96], mem[97], mem[98], mem[99], 
        mem[100], mem[101]}), .D3({mem[102], mem[103], mem[104], mem[105], 
        mem[106], mem[107], mem[108], mem[109], mem[110], mem[111], mem[112], 
        mem[113], mem[114], mem[115], mem[116], mem[117], mem[118], mem[119], 
        mem[120], mem[121], mem[122], mem[123], mem[124], mem[125], mem[126], 
        mem[127], mem[128], mem[129], mem[130], mem[131], mem[132], mem[133], 
        mem[134], mem[135]}), .D4({mem[136], mem[137], mem[138], mem[139], 
        mem[140], mem[141], mem[142], mem[143], mem[144], mem[145], mem[146], 
        mem[147], mem[148], mem[149], mem[150], mem[151], mem[152], mem[153], 
        mem[154], mem[155], mem[156], mem[157], mem[158], mem[159], mem[160], 
        mem[161], mem[162], mem[163], mem[164], mem[165], mem[166], mem[167], 
        mem[168], mem[169]}), .D5({mem[170], mem[171], mem[172], mem[173], 
        mem[174], mem[175], mem[176], mem[177], mem[178], mem[179], mem[180], 
        mem[181], mem[182], mem[183], mem[184], mem[185], mem[186], mem[187], 
        mem[188], mem[189], mem[190], mem[191], mem[192], mem[193], mem[194], 
        mem[195], mem[196], mem[197], mem[198], mem[199], mem[200], mem[201], 
        mem[202], mem[203]}), .D6({mem[204], mem[205], mem[206], mem[207], 
        mem[208], mem[209], mem[210], mem[211], mem[212], mem[213], mem[214], 
        mem[215], mem[216], mem[217], mem[218], mem[219], mem[220], mem[221], 
        mem[222], mem[223], mem[224], mem[225], mem[226], mem[227], mem[228], 
        mem[229], mem[230], mem[231], mem[232], mem[233], mem[234], mem[235], 
        mem[236], mem[237]}), .D7({mem[238], mem[239], mem[240], mem[241], 
        mem[242], mem[243], mem[244], mem[245], mem[246], mem[247], mem[248], 
        mem[249], mem[250], mem[251], mem[252], mem[253], mem[254], mem[255], 
        mem[256], mem[257], mem[258], mem[259], mem[260], mem[261], mem[262], 
        mem[263], mem[264], mem[265], mem[266], mem[267], mem[268], mem[269], 
        mem[270], mem[271]}), .D8({mem[272], mem[273], mem[274], mem[275], 
        mem[276], mem[277], mem[278], mem[279], mem[280], mem[281], mem[282], 
        mem[283], mem[284], mem[285], mem[286], mem[287], mem[288], mem[289], 
        mem[290], mem[291], mem[292], mem[293], mem[294], mem[295], mem[296], 
        mem[297], mem[298], mem[299], mem[300], mem[301], mem[302], mem[303], 
        mem[304], mem[305]}), .D9({mem[306], mem[307], mem[308], mem[309], 
        mem[310], mem[311], mem[312], mem[313], mem[314], mem[315], mem[316], 
        mem[317], mem[318], mem[319], mem[320], mem[321], mem[322], mem[323], 
        mem[324], mem[325], mem[326], mem[327], mem[328], mem[329], mem[330], 
        mem[331], mem[332], mem[333], mem[334], mem[335], mem[336], mem[337], 
        mem[338], mem[339]}), .D10({mem[340], mem[341], mem[342], mem[343], 
        mem[344], mem[345], mem[346], mem[347], mem[348], mem[349], mem[350], 
        mem[351], mem[352], mem[353], mem[354], mem[355], mem[356], mem[357], 
        mem[358], mem[359], mem[360], mem[361], mem[362], mem[363], mem[364], 
        mem[365], mem[366], mem[367], mem[368], mem[369], mem[370], mem[371], 
        mem[372], mem[373]}), .D11({mem[374], mem[375], mem[376], mem[377], 
        mem[378], mem[379], mem[380], mem[381], mem[382], mem[383], mem[384], 
        mem[385], mem[386], mem[387], mem[388], mem[389], mem[390], mem[391], 
        mem[392], mem[393], mem[394], mem[395], mem[396], mem[397], mem[398], 
        mem[399], mem[400], mem[401], mem[402], mem[403], mem[404], mem[405], 
        mem[406], mem[407]}), .D12({mem[408], mem[409], mem[410], mem[411], 
        mem[412], mem[413], mem[414], mem[415], mem[416], mem[417], mem[418], 
        mem[419], mem[420], mem[421], mem[422], mem[423], mem[424], mem[425], 
        mem[426], mem[427], mem[428], mem[429], mem[430], mem[431], mem[432], 
        mem[433], mem[434], mem[435], mem[436], mem[437], mem[438], mem[439], 
        mem[440], mem[441]}), .D13({mem[442], mem[443], mem[444], mem[445], 
        mem[446], mem[447], mem[448], mem[449], mem[450], mem[451], mem[452], 
        mem[453], mem[454], mem[455], mem[456], mem[457], mem[458], mem[459], 
        mem[460], mem[461], mem[462], mem[463], mem[464], mem[465], mem[466], 
        mem[467], mem[468], mem[469], mem[470], mem[471], mem[472], mem[473], 
        mem[474], mem[475]}), .D14({mem[476], mem[477], mem[478], mem[479], 
        mem[480], mem[481], mem[482], mem[483], mem[484], mem[485], mem[486], 
        mem[487], mem[488], mem[489], mem[490], mem[491], mem[492], mem[493], 
        mem[494], mem[495], mem[496], mem[497], mem[498], mem[499], mem[500], 
        mem[501], mem[502], mem[503], mem[504], mem[505], mem[506], mem[507], 
        mem[508], mem[509]}), .D15({mem[510], mem[511], mem[512], mem[513], 
        mem[514], mem[515], mem[516], mem[517], mem[518], mem[519], mem[520], 
        mem[521], mem[522], mem[523], mem[524], mem[525], mem[526], mem[527], 
        mem[528], mem[529], mem[530], mem[531], mem[532], mem[533], mem[534], 
        mem[535], mem[536], mem[537], mem[538], mem[539], mem[540], mem[541], 
        mem[542], mem[543]}), .D16({mem[544], mem[545], mem[546], mem[547], 
        mem[548], mem[549], mem[550], mem[551], mem[552], mem[553], mem[554], 
        mem[555], mem[556], mem[557], mem[558], mem[559], mem[560], mem[561], 
        mem[562], mem[563], mem[564], mem[565], mem[566], mem[567], mem[568], 
        mem[569], mem[570], mem[571], mem[572], mem[573], mem[574], mem[575], 
        mem[576], mem[577]}), .D17({mem[578], mem[579], mem[580], mem[581], 
        mem[582], mem[583], mem[584], mem[585], mem[586], mem[587], mem[588], 
        mem[589], mem[590], mem[591], mem[592], mem[593], mem[594], mem[595], 
        mem[596], mem[597], mem[598], mem[599], mem[600], mem[601], mem[602], 
        mem[603], mem[604], mem[605], mem[606], mem[607], mem[608], mem[609], 
        mem[610], mem[611]}), .D18({mem[612], mem[613], mem[614], mem[615], 
        mem[616], mem[617], mem[618], mem[619], mem[620], mem[621], mem[622], 
        mem[623], mem[624], mem[625], mem[626], mem[627], mem[628], mem[629], 
        mem[630], mem[631], mem[632], mem[633], mem[634], mem[635], mem[636], 
        mem[637], mem[638], mem[639], mem[640], mem[641], mem[642], mem[643], 
        mem[644], mem[645]}), .D19({mem[646], mem[647], mem[648], mem[649], 
        mem[650], mem[651], mem[652], mem[653], mem[654], mem[655], mem[656], 
        mem[657], mem[658], mem[659], mem[660], mem[661], mem[662], mem[663], 
        mem[664], mem[665], mem[666], mem[667], mem[668], mem[669], mem[670], 
        mem[671], mem[672], mem[673], mem[674], mem[675], mem[676], mem[677], 
        mem[678], mem[679]}), .D20({mem[680], mem[681], mem[682], mem[683], 
        mem[684], mem[685], mem[686], mem[687], mem[688], mem[689], mem[690], 
        mem[691], mem[692], mem[693], mem[694], mem[695], mem[696], mem[697], 
        mem[698], mem[699], mem[700], mem[701], mem[702], mem[703], mem[704], 
        mem[705], mem[706], mem[707], mem[708], mem[709], mem[710], mem[711], 
        mem[712], mem[713]}), .D21({mem[714], mem[715], mem[716], mem[717], 
        mem[718], mem[719], mem[720], mem[721], mem[722], mem[723], mem[724], 
        mem[725], mem[726], mem[727], mem[728], mem[729], mem[730], mem[731], 
        mem[732], mem[733], mem[734], mem[735], mem[736], mem[737], mem[738], 
        mem[739], mem[740], mem[741], mem[742], mem[743], mem[744], mem[745], 
        mem[746], mem[747]}), .D22({mem[748], mem[749], mem[750], mem[751], 
        mem[752], mem[753], mem[754], mem[755], mem[756], mem[757], mem[758], 
        mem[759], mem[760], mem[761], mem[762], mem[763], mem[764], mem[765], 
        mem[766], mem[767], mem[768], mem[769], mem[770], mem[771], mem[772], 
        mem[773], mem[774], mem[775], mem[776], mem[777], mem[778], mem[779], 
        mem[780], mem[781]}), .D23({mem[782], mem[783], mem[784], mem[785], 
        mem[786], mem[787], mem[788], mem[789], mem[790], mem[791], mem[792], 
        mem[793], mem[794], mem[795], mem[796], mem[797], mem[798], mem[799], 
        mem[800], mem[801], mem[802], mem[803], mem[804], mem[805], mem[806], 
        mem[807], mem[808], mem[809], mem[810], mem[811], mem[812], mem[813], 
        mem[814], mem[815]}), .D24({mem[816], mem[817], mem[818], mem[819], 
        mem[820], mem[821], mem[822], mem[823], mem[824], mem[825], mem[826], 
        mem[827], mem[828], mem[829], mem[830], mem[831], mem[832], mem[833], 
        mem[834], mem[835], mem[836], mem[837], mem[838], mem[839], mem[840], 
        mem[841], mem[842], mem[843], mem[844], mem[845], mem[846], mem[847], 
        mem[848], mem[849]}), .D25({mem[850], mem[851], mem[852], mem[853], 
        mem[854], mem[855], mem[856], mem[857], mem[858], mem[859], mem[860], 
        mem[861], mem[862], mem[863], mem[864], mem[865], mem[866], mem[867], 
        mem[868], mem[869], mem[870], mem[871], mem[872], mem[873], mem[874], 
        mem[875], mem[876], mem[877], mem[878], mem[879], mem[880], mem[881], 
        mem[882], mem[883]}), .D26({mem[884], mem[885], mem[886], mem[887], 
        mem[888], mem[889], mem[890], mem[891], mem[892], mem[893], mem[894], 
        mem[895], mem[896], mem[897], mem[898], mem[899], mem[900], mem[901], 
        mem[902], mem[903], mem[904], mem[905], mem[906], mem[907], mem[908], 
        mem[909], mem[910], mem[911], mem[912], mem[913], mem[914], mem[915], 
        mem[916], mem[917]}), .D27({mem[918], mem[919], mem[920], mem[921], 
        mem[922], mem[923], mem[924], mem[925], mem[926], mem[927], mem[928], 
        mem[929], mem[930], mem[931], mem[932], mem[933], mem[934], mem[935], 
        mem[936], mem[937], mem[938], mem[939], mem[940], mem[941], mem[942], 
        mem[943], mem[944], mem[945], mem[946], mem[947], mem[948], mem[949], 
        mem[950], mem[951]}), .D28({mem[952], mem[953], mem[954], mem[955], 
        mem[956], mem[957], mem[958], mem[959], mem[960], mem[961], mem[962], 
        mem[963], mem[964], mem[965], mem[966], mem[967], mem[968], mem[969], 
        mem[970], mem[971], mem[972], mem[973], mem[974], mem[975], mem[976], 
        mem[977], mem[978], mem[979], mem[980], mem[981], mem[982], mem[983], 
        mem[984], mem[985]}), .D29({mem[986], mem[987], mem[988], mem[989], 
        mem[990], mem[991], mem[992], mem[993], mem[994], mem[995], mem[996], 
        mem[997], mem[998], mem[999], mem[1000], mem[1001], mem[1002], 
        mem[1003], mem[1004], mem[1005], mem[1006], mem[1007], mem[1008], 
        mem[1009], mem[1010], mem[1011], mem[1012], mem[1013], mem[1014], 
        mem[1015], mem[1016], mem[1017], mem[1018], mem[1019]}), .D30({
        mem[1020], mem[1021], mem[1022], mem[1023], mem[1024], mem[1025], 
        mem[1026], mem[1027], mem[1028], mem[1029], mem[1030], mem[1031], 
        mem[1032], mem[1033], mem[1034], mem[1035], mem[1036], mem[1037], 
        mem[1038], mem[1039], mem[1040], mem[1041], mem[1042], mem[1043], 
        mem[1044], mem[1045], mem[1046], mem[1047], mem[1048], mem[1049], 
        mem[1050], mem[1051], mem[1052], mem[1053]}), .D31({mem[1054], 
        mem[1055], mem[1056], mem[1057], mem[1058], mem[1059], mem[1060], 
        mem[1061], mem[1062], mem[1063], mem[1064], mem[1065], mem[1066], 
        mem[1067], mem[1068], mem[1069], mem[1070], mem[1071], mem[1072], 
        mem[1073], mem[1074], mem[1075], mem[1076], mem[1077], mem[1078], 
        mem[1079], mem[1080], mem[1081], mem[1082], mem[1083], mem[1084], 
        mem[1085], mem[1086], mem[1087]}), .S0(N18), .S1(N19), .S2(N20), .S3(
        N21), .S4(N22), .Z({data_out[0], data_out[1], data_out[2], data_out[3], 
        data_out[4], data_out[5], data_out[6], data_out[7], data_out[8], 
        data_out[9], data_out[10], data_out[11], data_out[12], data_out[13], 
        data_out[14], data_out[15], data_out[16], data_out[17], data_out[18], 
        data_out[19], data_out[20], data_out[21], data_out[22], data_out[23], 
        data_out[24], data_out[25], data_out[26], data_out[27], data_out[28], 
        data_out[29], data_out[30], data_out[31], data_out[32], data_out[33]})
         );
  GTECH_BUF B_2 ( .A(rd_ptr[0]), .Z(N18) );
  GTECH_BUF B_3 ( .A(rd_ptr[1]), .Z(N19) );
  GTECH_BUF B_4 ( .A(rd_ptr[2]), .Z(N20) );
  GTECH_BUF B_5 ( .A(rd_ptr[3]), .Z(N21) );
  GTECH_BUF B_6 ( .A(rd_ptr[4]), .Z(N22) );
  GTECH_AND2 C9210 ( .A(N228), .B(put), .Z(N23) );
  GTECH_NOT I_18 ( .A(fillcount[5]), .Z(N228) );
  GTECH_AND2 C9213 ( .A(N229), .B(get), .Z(N24) );
  GTECH_AND2 C9214 ( .A(N23), .B(N128), .Z(N229) );
  GTECH_AND2 C9215 ( .A(N128), .B(get), .Z(N25) );
  GTECH_OR2 C9220 ( .A(N24), .B(reset), .Z(N26) );
  GTECH_OR2 C9221 ( .A(N23), .B(N26), .Z(N27) );
  GTECH_OR2 C9222 ( .A(N25), .B(N27), .Z(N28) );
  GTECH_NOT I_19 ( .A(N28), .Z(N29) );
  GTECH_BUF B_7 ( .A(N117), .Z(N30) );
  GTECH_BUF B_8 ( .A(N120), .Z(N41) );
  GTECH_BUF B_9 ( .A(N123), .Z(N53) );
  GTECH_NOT I_20 ( .A(reset), .Z(N116) );
  GTECH_AND2 C9292 ( .A(N24), .B(N116), .Z(N117) );
  GTECH_AND2 C9293 ( .A(N30), .B(N116), .Z(net342) );
  GTECH_NOT I_21 ( .A(N24), .Z(N118) );
  GTECH_AND2 C9295 ( .A(N116), .B(N118), .Z(N119) );
  GTECH_AND2 C9296 ( .A(N23), .B(N119), .Z(N120) );
  GTECH_AND2 C9297 ( .A(N41), .B(N119), .Z(net343) );
  GTECH_NOT I_22 ( .A(N23), .Z(N121) );
  GTECH_AND2 C9299 ( .A(N119), .B(N121), .Z(N122) );
  GTECH_AND2 C9300 ( .A(N25), .B(N122), .Z(N123) );
  GTECH_AND2 C9301 ( .A(N53), .B(N122), .Z(net344) );
endmodule


module FIFO_DEPTH_P25_WIDTH42 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [41:0] data_in;
  output [41:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, net421, net422,
         net423;
  wire   [4:0] wr_ptr;
  wire   [4:0] rd_ptr;
  wire   [1343:0] mem;
  tri   clk;
  tri   reset;
  tri   [41:0] data_in;
  tri   put;
  tri   [5:0] fillcount;
  assign full = fillcount[5];

  \**SEQGEN**  mem_reg_31__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1343]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1342]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1341]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1340]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1339]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1338]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1337]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1336]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1335]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1334]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1333]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1332]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1331]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1330]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1329]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1328]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1327]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1326]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1325]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1324]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1323]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1322]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1321]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1320]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1319]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1318]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1317]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1316]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1315]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1314]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1313]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1312]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1311]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1310]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1309]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1308]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1307]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1306]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1305]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1304]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1303]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_31__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1302]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N115) );
  \**SEQGEN**  mem_reg_30__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1301]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1300]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1299]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1298]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1297]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1296]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1295]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1294]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1293]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1292]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1291]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1290]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1289]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1288]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1287]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1286]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1285]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1284]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1283]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1282]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1281]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1280]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1279]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1278]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1277]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1276]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1275]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1274]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1273]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1272]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1271]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1270]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1269]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1268]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1267]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1266]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1265]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1264]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1263]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1262]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1261]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_30__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1260]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N114) );
  \**SEQGEN**  mem_reg_29__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1259]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1258]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1257]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1256]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_29__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N113) );
  \**SEQGEN**  mem_reg_28__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_28__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N112) );
  \**SEQGEN**  mem_reg_27__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_27__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N111) );
  \**SEQGEN**  mem_reg_26__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1099]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1098]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1097]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1096]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1095]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1094]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1093]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_26__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1092]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N110) );
  \**SEQGEN**  mem_reg_25__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1091]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1090]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1089]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1088]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1087]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1086]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1085]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1084]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1083]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1082]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1081]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1080]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1079]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1078]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1077]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1076]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1075]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1074]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1073]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1072]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1071]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1070]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1069]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1068]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1067]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1066]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1065]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1064]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1063]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1062]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1061]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1060]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1059]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1058]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1057]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1056]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1055]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1054]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1053]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1052]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1051]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_25__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1050]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N109) );
  \**SEQGEN**  mem_reg_24__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1049]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1048]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1047]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1046]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1045]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1044]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1043]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1042]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1041]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1040]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1039]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1038]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1037]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1036]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1035]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1034]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1033]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1032]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1031]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1030]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1029]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1028]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1027]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1026]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1025]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1024]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1023]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1022]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1021]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1020]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1019]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1018]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1017]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1016]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1015]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1014]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1013]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1012]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1011]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1010]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1009]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_24__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1008]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N108) );
  \**SEQGEN**  mem_reg_23__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1007]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1006]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1005]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1004]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1003]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1002]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1001]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1000]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[999]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[998]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[997]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[996]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[995]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[994]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[993]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[992]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[991]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[990]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[989]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[988]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[987]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[986]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[985]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[984]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[983]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[982]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[981]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[980]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[979]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[978]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[977]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[976]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[975]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[974]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[973]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[972]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[971]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[970]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[969]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[968]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[967]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_23__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[966]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N107) );
  \**SEQGEN**  mem_reg_22__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[965]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[964]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[963]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[962]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[961]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[960]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[959]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[958]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[957]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[956]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[955]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[954]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[953]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[952]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[951]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[950]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[949]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[948]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[947]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[946]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[945]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[944]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[943]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[942]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[941]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[940]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[939]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[938]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[937]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[936]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[935]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[934]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[933]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[932]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[931]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[930]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[929]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[928]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[927]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[926]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[925]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_22__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[924]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N106) );
  \**SEQGEN**  mem_reg_21__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[923]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[922]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[921]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[920]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[919]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[918]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[917]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[916]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[915]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[914]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[913]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[912]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[911]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[910]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[909]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[908]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[907]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[906]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[905]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[904]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[903]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[902]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[901]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[900]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[899]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[898]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[897]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[896]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[895]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[894]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[893]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[892]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[891]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[890]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[889]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[888]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[887]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[886]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[885]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[884]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[883]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_21__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[882]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N105) );
  \**SEQGEN**  mem_reg_20__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[881]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[880]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[879]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[878]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[877]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[876]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[875]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[874]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[873]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[872]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[871]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[870]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[869]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[868]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[867]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[866]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[865]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[864]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[863]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[862]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[861]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[860]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[859]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[858]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[857]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[856]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[855]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[854]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[853]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[852]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[851]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[850]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[849]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[848]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[847]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[846]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[845]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[844]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[843]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[842]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[841]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_20__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[840]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N104) );
  \**SEQGEN**  mem_reg_19__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[839]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[838]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[837]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[836]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[835]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[834]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[833]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[832]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[831]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[830]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[829]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[828]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[827]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[826]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[825]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[824]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[823]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[822]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[821]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[820]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[819]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[818]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[817]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[816]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[815]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[814]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[813]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[812]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[811]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[810]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[809]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[808]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[807]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[806]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[805]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[804]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[803]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[802]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[801]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[800]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[799]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_19__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[798]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  mem_reg_18__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[797]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[796]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[795]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[794]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[793]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[792]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[791]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[790]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[789]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[788]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[787]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[786]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[785]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[784]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[783]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[782]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[781]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[780]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[779]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[778]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[777]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[776]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[775]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[774]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[773]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[772]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[771]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[770]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[769]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[768]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[767]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[766]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[765]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[764]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[763]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[762]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[761]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[760]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[759]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[758]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[757]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_18__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[756]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N102) );
  \**SEQGEN**  mem_reg_17__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[755]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[754]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[753]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[752]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[751]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[750]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[749]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[748]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[747]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[746]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[745]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[744]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[743]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[742]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[741]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[740]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[739]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[738]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[737]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[736]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[735]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[734]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[733]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[732]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[731]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[730]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[729]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[728]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[727]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[726]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[725]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[724]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[723]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[722]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[721]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[720]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[719]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[718]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[717]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[716]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[715]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_17__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[714]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N101) );
  \**SEQGEN**  mem_reg_16__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[713]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[712]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[711]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[710]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[709]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[708]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[707]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[706]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[705]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[704]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[703]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[702]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[701]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[700]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[699]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[698]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[697]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[696]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[695]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[694]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[693]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[692]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[691]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[690]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[689]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[688]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[687]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[686]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[685]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[684]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[683]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[682]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[681]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[680]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[679]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[678]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[677]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[676]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[675]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[674]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[673]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_16__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[672]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N100) );
  \**SEQGEN**  mem_reg_15__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[671]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[670]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[669]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[668]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[667]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[666]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[665]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[664]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[663]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[662]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[661]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[660]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[659]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[658]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[657]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[656]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[655]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[654]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[653]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[652]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[651]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[650]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[649]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[648]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[647]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[646]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[645]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[644]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[643]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[642]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[641]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[640]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[639]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[638]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[637]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[636]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[635]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[634]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[633]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[632]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[631]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_15__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[630]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N99) );
  \**SEQGEN**  mem_reg_14__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[629]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[628]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[627]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[626]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[625]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[624]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[623]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[622]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[621]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[620]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[619]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[618]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[617]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[616]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[615]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[614]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[613]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[612]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[611]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[610]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[609]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[608]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[607]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[606]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[605]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[604]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[603]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[602]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[601]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[600]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[599]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[598]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[597]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[596]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[595]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[594]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[593]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[592]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[591]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[590]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[589]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_14__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[588]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N98) );
  \**SEQGEN**  mem_reg_13__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[587]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[586]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[585]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[584]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[583]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[582]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[581]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[580]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[579]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[578]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[577]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[576]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[575]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[574]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[573]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[572]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[571]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[570]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[569]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[568]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[567]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[566]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[565]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[564]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[563]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[562]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[561]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[560]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[559]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[558]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[557]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[556]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[555]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[554]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[553]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[552]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[551]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[550]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[549]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[548]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[547]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_13__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[546]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N97) );
  \**SEQGEN**  mem_reg_12__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[545]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[544]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[543]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[542]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[541]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[540]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[539]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[538]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[537]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[536]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[535]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[534]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[533]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[532]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[531]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[530]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[529]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[528]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[527]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[526]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[525]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[524]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[523]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[522]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[521]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[520]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[519]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[518]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[517]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[516]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[515]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[514]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[513]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[512]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[511]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[510]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[509]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[508]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[507]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[506]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[505]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_12__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[504]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N96) );
  \**SEQGEN**  mem_reg_11__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[503]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[502]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[501]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[500]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[499]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[498]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[497]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[496]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[495]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[494]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[493]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[492]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[491]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[490]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[489]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[488]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[487]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[486]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[485]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[484]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[483]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[482]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[481]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[480]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[479]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[478]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[477]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[476]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[475]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[474]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[473]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[472]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[471]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[470]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[469]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[468]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[467]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[466]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[465]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[464]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[463]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_11__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[462]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N95) );
  \**SEQGEN**  mem_reg_10__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[461]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[460]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[459]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[458]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[457]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[456]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[455]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[454]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[453]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[452]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[451]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[450]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[449]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[448]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[447]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[446]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[445]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[444]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[443]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[442]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[441]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[440]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[439]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[438]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[437]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[436]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[435]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[434]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[433]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[432]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[431]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[430]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[429]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[428]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[427]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[426]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[425]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[424]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[423]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[422]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[421]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_10__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[420]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N94) );
  \**SEQGEN**  mem_reg_9__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[419]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[418]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[417]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[416]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[415]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[414]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[413]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[412]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[411]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[410]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[409]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[408]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[407]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[406]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[405]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[404]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[403]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[402]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[401]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[400]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[399]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[398]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[397]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[396]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[395]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[394]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[393]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[392]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[391]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[390]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[389]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[388]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[387]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[386]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[385]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[384]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[383]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[382]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[381]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[380]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[379]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_9__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[378]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N93) );
  \**SEQGEN**  mem_reg_8__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[377]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[376]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[375]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[374]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[373]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[372]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[371]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[370]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[369]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[368]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[367]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[366]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[365]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[364]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[363]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[362]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[361]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[360]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[359]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[358]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[357]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[356]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[355]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[354]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[353]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[352]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[351]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[350]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[349]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[348]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[347]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[346]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[345]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[344]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[343]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[342]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[341]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[340]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[339]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[338]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[337]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_8__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[336]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N92) );
  \**SEQGEN**  mem_reg_7__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[335]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[334]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[333]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[332]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[331]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[330]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[329]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[328]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[327]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[326]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[325]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[324]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[323]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[322]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[321]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[320]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[319]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[318]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[317]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[316]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[315]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[314]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[313]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[312]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[311]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[310]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[309]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[308]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[307]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[306]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[305]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[304]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[303]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[302]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[301]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[300]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[299]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[298]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[297]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[296]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[295]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_7__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[294]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N91) );
  \**SEQGEN**  mem_reg_6__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[293]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[292]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[291]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[290]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[289]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[288]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[287]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[286]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[285]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[284]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[283]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[282]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[281]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[280]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[279]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[278]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[277]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[276]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[275]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[274]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[273]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[272]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[271]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[270]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[269]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[268]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[267]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[266]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[265]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[264]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[263]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[262]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[261]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[260]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[259]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[258]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[257]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[256]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_6__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N90) );
  \**SEQGEN**  mem_reg_5__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_5__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N89) );
  \**SEQGEN**  mem_reg_4__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_4__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N88) );
  \**SEQGEN**  mem_reg_3__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_3__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N87) );
  \**SEQGEN**  mem_reg_2__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[99]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[98]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[97]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[96]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[95]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[94]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[93]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[92]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[91]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[90]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[89]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[88]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[87]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[86]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[85]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_2__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[84]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N86) );
  \**SEQGEN**  mem_reg_1__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[83]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[82]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[81]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[80]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[79]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[78]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[77]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[76]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[75]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[74]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[73]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[72]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[71]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[70]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[69]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[68]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[67]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[66]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[65]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[64]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[63]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[62]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[61]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[60]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[59]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[58]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[57]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[56]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[55]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[54]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[53]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[52]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[51]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[50]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[49]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[48]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[47]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[46]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[45]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[44]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[43]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_1__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[42]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N85) );
  \**SEQGEN**  mem_reg_0__41_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[41]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__40_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[40]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__39_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[39]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__38_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[38]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__37_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[37]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__36_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[36]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__35_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[35]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__34_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[34]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__33_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[33]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__32_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[32]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__31_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__30_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__29_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__28_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__27_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__26_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__25_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__24_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__23_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__22_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__21_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__20_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__19_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__18_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__17_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__16_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__15_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__14_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__13_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__12_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__11_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__9_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__8_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  mem_reg_0__0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        data_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        mem[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N84) );
  \**SEQGEN**  fillcount_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N83), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N82), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N81), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N80), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N79), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  fillcount_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N78), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(fillcount[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N77) );
  \**SEQGEN**  rd_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  rd_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rd_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  wr_ptr_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  \**SEQGEN**  wr_ptr_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(wr_ptr[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N65) );
  GTECH_OR2 C8411 ( .A(fillcount[4]), .B(fillcount[5]), .Z(N124) );
  GTECH_OR2 C8412 ( .A(fillcount[3]), .B(N124), .Z(N125) );
  GTECH_OR2 C8413 ( .A(fillcount[2]), .B(N125), .Z(N126) );
  GTECH_OR2 C8414 ( .A(fillcount[1]), .B(N126), .Z(N127) );
  GTECH_OR2 C8415 ( .A(fillcount[0]), .B(N127), .Z(N128) );
  GTECH_NOT I_0 ( .A(N128), .Z(empty) );
  ADD_UNS_OP add_33 ( .A(rd_ptr), .B(1'b1), .Z({N40, N39, N38, N37, N36}) );
  ADD_UNS_OP add_32 ( .A(wr_ptr), .B(1'b1), .Z({N35, N34, N33, N32, N31}) );
  GTECH_OR3 C8417 ( .A(reset), .B(N117), .C(N120), .Z(N65) );
  GTECH_OR3 C8432 ( .A(reset), .B(N117), .C(N123), .Z(N71) );
  GTECH_OR3 C8447 ( .A(reset), .B(N120), .C(N123), .Z(N77) );
  ADD_UNS_OP add_37 ( .A(fillcount), .B(1'b1), .Z({N52, N51, N50, N49, N48, 
        N47}) );
  ADD_UNS_OP add_36 ( .A(wr_ptr), .B(1'b1), .Z({N46, N45, N44, N43, N42}) );
  SUB_UNS_OP sub_40 ( .A(fillcount), .B(1'b1), .Z({N64, N63, N62, N61, N60, 
        N59}) );
  ADD_UNS_OP add_39 ( .A(rd_ptr), .B(1'b1), .Z({N58, N57, N56, N55, N54}) );
  GTECH_OR3 C8465 ( .A(reset), .B(N123), .C(N29), .Z(N130) );
  GTECH_AND2 C11153 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N131) );
  GTECH_AND2 C11154 ( .A(N0), .B(wr_ptr[4]), .Z(N132) );
  GTECH_NOT I_1 ( .A(wr_ptr[3]), .Z(N0) );
  GTECH_AND2 C11155 ( .A(wr_ptr[3]), .B(N1), .Z(N133) );
  GTECH_NOT I_2 ( .A(wr_ptr[4]), .Z(N1) );
  GTECH_AND2 C11156 ( .A(N2), .B(N3), .Z(N134) );
  GTECH_NOT I_3 ( .A(wr_ptr[3]), .Z(N2) );
  GTECH_NOT I_4 ( .A(wr_ptr[4]), .Z(N3) );
  GTECH_NOT I_5 ( .A(wr_ptr[2]), .Z(N135) );
  GTECH_AND2 C11158 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N136) );
  GTECH_AND2 C11159 ( .A(N4), .B(wr_ptr[1]), .Z(N137) );
  GTECH_NOT I_6 ( .A(wr_ptr[0]), .Z(N4) );
  GTECH_AND2 C11160 ( .A(wr_ptr[0]), .B(N5), .Z(N138) );
  GTECH_NOT I_7 ( .A(wr_ptr[1]), .Z(N5) );
  GTECH_AND2 C11161 ( .A(N6), .B(N7), .Z(N139) );
  GTECH_NOT I_8 ( .A(wr_ptr[0]), .Z(N6) );
  GTECH_NOT I_9 ( .A(wr_ptr[1]), .Z(N7) );
  GTECH_AND2 C11162 ( .A(wr_ptr[2]), .B(N136), .Z(N140) );
  GTECH_AND2 C11163 ( .A(wr_ptr[2]), .B(N137), .Z(N141) );
  GTECH_AND2 C11164 ( .A(wr_ptr[2]), .B(N138), .Z(N142) );
  GTECH_AND2 C11165 ( .A(wr_ptr[2]), .B(N139), .Z(N143) );
  GTECH_AND2 C11166 ( .A(N135), .B(N136), .Z(N144) );
  GTECH_AND2 C11167 ( .A(N135), .B(N137), .Z(N145) );
  GTECH_AND2 C11168 ( .A(N135), .B(N138), .Z(N146) );
  GTECH_AND2 C11169 ( .A(N135), .B(N139), .Z(N147) );
  GTECH_AND2 C11170 ( .A(N131), .B(N140), .Z(N148) );
  GTECH_AND2 C11171 ( .A(N131), .B(N141), .Z(N149) );
  GTECH_AND2 C11172 ( .A(N131), .B(N142), .Z(N150) );
  GTECH_AND2 C11173 ( .A(N131), .B(N143), .Z(N151) );
  GTECH_AND2 C11174 ( .A(N131), .B(N144), .Z(N152) );
  GTECH_AND2 C11175 ( .A(N131), .B(N145), .Z(N153) );
  GTECH_AND2 C11176 ( .A(N131), .B(N146), .Z(N154) );
  GTECH_AND2 C11177 ( .A(N131), .B(N147), .Z(N155) );
  GTECH_AND2 C11178 ( .A(N132), .B(N140), .Z(N156) );
  GTECH_AND2 C11179 ( .A(N132), .B(N141), .Z(N157) );
  GTECH_AND2 C11180 ( .A(N132), .B(N142), .Z(N158) );
  GTECH_AND2 C11181 ( .A(N132), .B(N143), .Z(N159) );
  GTECH_AND2 C11182 ( .A(N132), .B(N144), .Z(N160) );
  GTECH_AND2 C11183 ( .A(N132), .B(N145), .Z(N161) );
  GTECH_AND2 C11184 ( .A(N132), .B(N146), .Z(N162) );
  GTECH_AND2 C11185 ( .A(N132), .B(N147), .Z(N163) );
  GTECH_AND2 C11186 ( .A(N133), .B(N140), .Z(N164) );
  GTECH_AND2 C11187 ( .A(N133), .B(N141), .Z(N165) );
  GTECH_AND2 C11188 ( .A(N133), .B(N142), .Z(N166) );
  GTECH_AND2 C11189 ( .A(N133), .B(N143), .Z(N167) );
  GTECH_AND2 C11190 ( .A(N133), .B(N144), .Z(N168) );
  GTECH_AND2 C11191 ( .A(N133), .B(N145), .Z(N169) );
  GTECH_AND2 C11192 ( .A(N133), .B(N146), .Z(N170) );
  GTECH_AND2 C11193 ( .A(N133), .B(N147), .Z(N171) );
  GTECH_AND2 C11194 ( .A(N134), .B(N140), .Z(N172) );
  GTECH_AND2 C11195 ( .A(N134), .B(N141), .Z(N173) );
  GTECH_AND2 C11196 ( .A(N134), .B(N142), .Z(N174) );
  GTECH_AND2 C11197 ( .A(N134), .B(N143), .Z(N175) );
  GTECH_AND2 C11198 ( .A(N134), .B(N144), .Z(N176) );
  GTECH_AND2 C11199 ( .A(N134), .B(N145), .Z(N177) );
  GTECH_AND2 C11200 ( .A(N134), .B(N146), .Z(N178) );
  GTECH_AND2 C11201 ( .A(N134), .B(N147), .Z(N179) );
  GTECH_AND2 C11202 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Z(N180) );
  GTECH_AND2 C11203 ( .A(N8), .B(wr_ptr[4]), .Z(N181) );
  GTECH_NOT I_10 ( .A(wr_ptr[3]), .Z(N8) );
  GTECH_AND2 C11204 ( .A(wr_ptr[3]), .B(N9), .Z(N182) );
  GTECH_NOT I_11 ( .A(wr_ptr[4]), .Z(N9) );
  GTECH_AND2 C11205 ( .A(N10), .B(N11), .Z(N183) );
  GTECH_NOT I_12 ( .A(wr_ptr[3]), .Z(N10) );
  GTECH_NOT I_13 ( .A(wr_ptr[4]), .Z(N11) );
  GTECH_AND2 C11207 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Z(N184) );
  GTECH_AND2 C11208 ( .A(N12), .B(wr_ptr[1]), .Z(N185) );
  GTECH_NOT I_14 ( .A(wr_ptr[0]), .Z(N12) );
  GTECH_AND2 C11209 ( .A(wr_ptr[0]), .B(N13), .Z(N186) );
  GTECH_NOT I_15 ( .A(wr_ptr[1]), .Z(N13) );
  GTECH_AND2 C11210 ( .A(N14), .B(N15), .Z(N187) );
  GTECH_NOT I_16 ( .A(wr_ptr[0]), .Z(N14) );
  GTECH_NOT I_17 ( .A(wr_ptr[1]), .Z(N15) );
  GTECH_AND2 C11211 ( .A(wr_ptr[2]), .B(N184), .Z(N188) );
  GTECH_AND2 C11212 ( .A(wr_ptr[2]), .B(N185), .Z(N189) );
  GTECH_AND2 C11213 ( .A(wr_ptr[2]), .B(N186), .Z(N190) );
  GTECH_AND2 C11214 ( .A(wr_ptr[2]), .B(N187), .Z(N191) );
  GTECH_AND2 C11215 ( .A(N135), .B(N184), .Z(N192) );
  GTECH_AND2 C11216 ( .A(N135), .B(N185), .Z(N193) );
  GTECH_AND2 C11217 ( .A(N135), .B(N186), .Z(N194) );
  GTECH_AND2 C11218 ( .A(N135), .B(N187), .Z(N195) );
  GTECH_AND2 C11219 ( .A(N180), .B(N188), .Z(N196) );
  GTECH_AND2 C11220 ( .A(N180), .B(N189), .Z(N197) );
  GTECH_AND2 C11221 ( .A(N180), .B(N190), .Z(N198) );
  GTECH_AND2 C11222 ( .A(N180), .B(N191), .Z(N199) );
  GTECH_AND2 C11223 ( .A(N180), .B(N192), .Z(N200) );
  GTECH_AND2 C11224 ( .A(N180), .B(N193), .Z(N201) );
  GTECH_AND2 C11225 ( .A(N180), .B(N194), .Z(N202) );
  GTECH_AND2 C11226 ( .A(N180), .B(N195), .Z(N203) );
  GTECH_AND2 C11227 ( .A(N181), .B(N188), .Z(N204) );
  GTECH_AND2 C11228 ( .A(N181), .B(N189), .Z(N205) );
  GTECH_AND2 C11229 ( .A(N181), .B(N190), .Z(N206) );
  GTECH_AND2 C11230 ( .A(N181), .B(N191), .Z(N207) );
  GTECH_AND2 C11231 ( .A(N181), .B(N192), .Z(N208) );
  GTECH_AND2 C11232 ( .A(N181), .B(N193), .Z(N209) );
  GTECH_AND2 C11233 ( .A(N181), .B(N194), .Z(N210) );
  GTECH_AND2 C11234 ( .A(N181), .B(N195), .Z(N211) );
  GTECH_AND2 C11235 ( .A(N182), .B(N188), .Z(N212) );
  GTECH_AND2 C11236 ( .A(N182), .B(N189), .Z(N213) );
  GTECH_AND2 C11237 ( .A(N182), .B(N190), .Z(N214) );
  GTECH_AND2 C11238 ( .A(N182), .B(N191), .Z(N215) );
  GTECH_AND2 C11239 ( .A(N182), .B(N192), .Z(N216) );
  GTECH_AND2 C11240 ( .A(N182), .B(N193), .Z(N217) );
  GTECH_AND2 C11241 ( .A(N182), .B(N194), .Z(N218) );
  GTECH_AND2 C11242 ( .A(N182), .B(N195), .Z(N219) );
  GTECH_AND2 C11243 ( .A(N183), .B(N188), .Z(N220) );
  GTECH_AND2 C11244 ( .A(N183), .B(N189), .Z(N221) );
  GTECH_AND2 C11245 ( .A(N183), .B(N190), .Z(N222) );
  GTECH_AND2 C11246 ( .A(N183), .B(N191), .Z(N223) );
  GTECH_AND2 C11247 ( .A(N183), .B(N192), .Z(N224) );
  GTECH_AND2 C11248 ( .A(N183), .B(N193), .Z(N225) );
  GTECH_AND2 C11249 ( .A(N183), .B(N194), .Z(N226) );
  GTECH_AND2 C11250 ( .A(N183), .B(N195), .Z(N227) );
  SELECT_OP C11251 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N35, N34, 
        N33, N32, N31}), .DATA3({N46, N45, N44, N43, N42}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N120), .Z({N70, N69, N68, N67, N66}) );
  GTECH_BUF B_0 ( .A(reset), .Z(N16) );
  SELECT_OP C11252 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N40, N39, 
        N38, N37, N36}), .DATA3({N58, N57, N56, N55, N54}), .CONTROL1(N16), 
        .CONTROL2(N117), .CONTROL3(N123), .Z({N76, N75, N74, N73, N72}) );
  SELECT_OP C11253 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N52, 
        N51, N50, N49, N48, N47}), .DATA3({N64, N63, N62, N61, N60, N59}), 
        .CONTROL1(N16), .CONTROL2(N120), .CONTROL3(N123), .Z({N83, N82, N81, 
        N80, N79, N78}) );
  SELECT_OP C11254 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
        N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
        N171, N172, N173, N174, N175, N176, N177, N178, N179}), .DATA3({N196, 
        N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
        N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
        N221, N222, N223, N224, N225, N226, N227}), .CONTROL1(N17), .CONTROL2(
        N117), .CONTROL3(N120), .Z({N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84}) );
  GTECH_BUF B_1 ( .A(N130), .Z(N17) );
  MUX_OP C11255 ( .D0({mem[0], mem[1], mem[2], mem[3], mem[4], mem[5], mem[6], 
        mem[7], mem[8], mem[9], mem[10], mem[11], mem[12], mem[13], mem[14], 
        mem[15], mem[16], mem[17], mem[18], mem[19], mem[20], mem[21], mem[22], 
        mem[23], mem[24], mem[25], mem[26], mem[27], mem[28], mem[29], mem[30], 
        mem[31], mem[32], mem[33], mem[34], mem[35], mem[36], mem[37], mem[38], 
        mem[39], mem[40], mem[41]}), .D1({mem[42], mem[43], mem[44], mem[45], 
        mem[46], mem[47], mem[48], mem[49], mem[50], mem[51], mem[52], mem[53], 
        mem[54], mem[55], mem[56], mem[57], mem[58], mem[59], mem[60], mem[61], 
        mem[62], mem[63], mem[64], mem[65], mem[66], mem[67], mem[68], mem[69], 
        mem[70], mem[71], mem[72], mem[73], mem[74], mem[75], mem[76], mem[77], 
        mem[78], mem[79], mem[80], mem[81], mem[82], mem[83]}), .D2({mem[84], 
        mem[85], mem[86], mem[87], mem[88], mem[89], mem[90], mem[91], mem[92], 
        mem[93], mem[94], mem[95], mem[96], mem[97], mem[98], mem[99], 
        mem[100], mem[101], mem[102], mem[103], mem[104], mem[105], mem[106], 
        mem[107], mem[108], mem[109], mem[110], mem[111], mem[112], mem[113], 
        mem[114], mem[115], mem[116], mem[117], mem[118], mem[119], mem[120], 
        mem[121], mem[122], mem[123], mem[124], mem[125]}), .D3({mem[126], 
        mem[127], mem[128], mem[129], mem[130], mem[131], mem[132], mem[133], 
        mem[134], mem[135], mem[136], mem[137], mem[138], mem[139], mem[140], 
        mem[141], mem[142], mem[143], mem[144], mem[145], mem[146], mem[147], 
        mem[148], mem[149], mem[150], mem[151], mem[152], mem[153], mem[154], 
        mem[155], mem[156], mem[157], mem[158], mem[159], mem[160], mem[161], 
        mem[162], mem[163], mem[164], mem[165], mem[166], mem[167]}), .D4({
        mem[168], mem[169], mem[170], mem[171], mem[172], mem[173], mem[174], 
        mem[175], mem[176], mem[177], mem[178], mem[179], mem[180], mem[181], 
        mem[182], mem[183], mem[184], mem[185], mem[186], mem[187], mem[188], 
        mem[189], mem[190], mem[191], mem[192], mem[193], mem[194], mem[195], 
        mem[196], mem[197], mem[198], mem[199], mem[200], mem[201], mem[202], 
        mem[203], mem[204], mem[205], mem[206], mem[207], mem[208], mem[209]}), 
        .D5({mem[210], mem[211], mem[212], mem[213], mem[214], mem[215], 
        mem[216], mem[217], mem[218], mem[219], mem[220], mem[221], mem[222], 
        mem[223], mem[224], mem[225], mem[226], mem[227], mem[228], mem[229], 
        mem[230], mem[231], mem[232], mem[233], mem[234], mem[235], mem[236], 
        mem[237], mem[238], mem[239], mem[240], mem[241], mem[242], mem[243], 
        mem[244], mem[245], mem[246], mem[247], mem[248], mem[249], mem[250], 
        mem[251]}), .D6({mem[252], mem[253], mem[254], mem[255], mem[256], 
        mem[257], mem[258], mem[259], mem[260], mem[261], mem[262], mem[263], 
        mem[264], mem[265], mem[266], mem[267], mem[268], mem[269], mem[270], 
        mem[271], mem[272], mem[273], mem[274], mem[275], mem[276], mem[277], 
        mem[278], mem[279], mem[280], mem[281], mem[282], mem[283], mem[284], 
        mem[285], mem[286], mem[287], mem[288], mem[289], mem[290], mem[291], 
        mem[292], mem[293]}), .D7({mem[294], mem[295], mem[296], mem[297], 
        mem[298], mem[299], mem[300], mem[301], mem[302], mem[303], mem[304], 
        mem[305], mem[306], mem[307], mem[308], mem[309], mem[310], mem[311], 
        mem[312], mem[313], mem[314], mem[315], mem[316], mem[317], mem[318], 
        mem[319], mem[320], mem[321], mem[322], mem[323], mem[324], mem[325], 
        mem[326], mem[327], mem[328], mem[329], mem[330], mem[331], mem[332], 
        mem[333], mem[334], mem[335]}), .D8({mem[336], mem[337], mem[338], 
        mem[339], mem[340], mem[341], mem[342], mem[343], mem[344], mem[345], 
        mem[346], mem[347], mem[348], mem[349], mem[350], mem[351], mem[352], 
        mem[353], mem[354], mem[355], mem[356], mem[357], mem[358], mem[359], 
        mem[360], mem[361], mem[362], mem[363], mem[364], mem[365], mem[366], 
        mem[367], mem[368], mem[369], mem[370], mem[371], mem[372], mem[373], 
        mem[374], mem[375], mem[376], mem[377]}), .D9({mem[378], mem[379], 
        mem[380], mem[381], mem[382], mem[383], mem[384], mem[385], mem[386], 
        mem[387], mem[388], mem[389], mem[390], mem[391], mem[392], mem[393], 
        mem[394], mem[395], mem[396], mem[397], mem[398], mem[399], mem[400], 
        mem[401], mem[402], mem[403], mem[404], mem[405], mem[406], mem[407], 
        mem[408], mem[409], mem[410], mem[411], mem[412], mem[413], mem[414], 
        mem[415], mem[416], mem[417], mem[418], mem[419]}), .D10({mem[420], 
        mem[421], mem[422], mem[423], mem[424], mem[425], mem[426], mem[427], 
        mem[428], mem[429], mem[430], mem[431], mem[432], mem[433], mem[434], 
        mem[435], mem[436], mem[437], mem[438], mem[439], mem[440], mem[441], 
        mem[442], mem[443], mem[444], mem[445], mem[446], mem[447], mem[448], 
        mem[449], mem[450], mem[451], mem[452], mem[453], mem[454], mem[455], 
        mem[456], mem[457], mem[458], mem[459], mem[460], mem[461]}), .D11({
        mem[462], mem[463], mem[464], mem[465], mem[466], mem[467], mem[468], 
        mem[469], mem[470], mem[471], mem[472], mem[473], mem[474], mem[475], 
        mem[476], mem[477], mem[478], mem[479], mem[480], mem[481], mem[482], 
        mem[483], mem[484], mem[485], mem[486], mem[487], mem[488], mem[489], 
        mem[490], mem[491], mem[492], mem[493], mem[494], mem[495], mem[496], 
        mem[497], mem[498], mem[499], mem[500], mem[501], mem[502], mem[503]}), 
        .D12({mem[504], mem[505], mem[506], mem[507], mem[508], mem[509], 
        mem[510], mem[511], mem[512], mem[513], mem[514], mem[515], mem[516], 
        mem[517], mem[518], mem[519], mem[520], mem[521], mem[522], mem[523], 
        mem[524], mem[525], mem[526], mem[527], mem[528], mem[529], mem[530], 
        mem[531], mem[532], mem[533], mem[534], mem[535], mem[536], mem[537], 
        mem[538], mem[539], mem[540], mem[541], mem[542], mem[543], mem[544], 
        mem[545]}), .D13({mem[546], mem[547], mem[548], mem[549], mem[550], 
        mem[551], mem[552], mem[553], mem[554], mem[555], mem[556], mem[557], 
        mem[558], mem[559], mem[560], mem[561], mem[562], mem[563], mem[564], 
        mem[565], mem[566], mem[567], mem[568], mem[569], mem[570], mem[571], 
        mem[572], mem[573], mem[574], mem[575], mem[576], mem[577], mem[578], 
        mem[579], mem[580], mem[581], mem[582], mem[583], mem[584], mem[585], 
        mem[586], mem[587]}), .D14({mem[588], mem[589], mem[590], mem[591], 
        mem[592], mem[593], mem[594], mem[595], mem[596], mem[597], mem[598], 
        mem[599], mem[600], mem[601], mem[602], mem[603], mem[604], mem[605], 
        mem[606], mem[607], mem[608], mem[609], mem[610], mem[611], mem[612], 
        mem[613], mem[614], mem[615], mem[616], mem[617], mem[618], mem[619], 
        mem[620], mem[621], mem[622], mem[623], mem[624], mem[625], mem[626], 
        mem[627], mem[628], mem[629]}), .D15({mem[630], mem[631], mem[632], 
        mem[633], mem[634], mem[635], mem[636], mem[637], mem[638], mem[639], 
        mem[640], mem[641], mem[642], mem[643], mem[644], mem[645], mem[646], 
        mem[647], mem[648], mem[649], mem[650], mem[651], mem[652], mem[653], 
        mem[654], mem[655], mem[656], mem[657], mem[658], mem[659], mem[660], 
        mem[661], mem[662], mem[663], mem[664], mem[665], mem[666], mem[667], 
        mem[668], mem[669], mem[670], mem[671]}), .D16({mem[672], mem[673], 
        mem[674], mem[675], mem[676], mem[677], mem[678], mem[679], mem[680], 
        mem[681], mem[682], mem[683], mem[684], mem[685], mem[686], mem[687], 
        mem[688], mem[689], mem[690], mem[691], mem[692], mem[693], mem[694], 
        mem[695], mem[696], mem[697], mem[698], mem[699], mem[700], mem[701], 
        mem[702], mem[703], mem[704], mem[705], mem[706], mem[707], mem[708], 
        mem[709], mem[710], mem[711], mem[712], mem[713]}), .D17({mem[714], 
        mem[715], mem[716], mem[717], mem[718], mem[719], mem[720], mem[721], 
        mem[722], mem[723], mem[724], mem[725], mem[726], mem[727], mem[728], 
        mem[729], mem[730], mem[731], mem[732], mem[733], mem[734], mem[735], 
        mem[736], mem[737], mem[738], mem[739], mem[740], mem[741], mem[742], 
        mem[743], mem[744], mem[745], mem[746], mem[747], mem[748], mem[749], 
        mem[750], mem[751], mem[752], mem[753], mem[754], mem[755]}), .D18({
        mem[756], mem[757], mem[758], mem[759], mem[760], mem[761], mem[762], 
        mem[763], mem[764], mem[765], mem[766], mem[767], mem[768], mem[769], 
        mem[770], mem[771], mem[772], mem[773], mem[774], mem[775], mem[776], 
        mem[777], mem[778], mem[779], mem[780], mem[781], mem[782], mem[783], 
        mem[784], mem[785], mem[786], mem[787], mem[788], mem[789], mem[790], 
        mem[791], mem[792], mem[793], mem[794], mem[795], mem[796], mem[797]}), 
        .D19({mem[798], mem[799], mem[800], mem[801], mem[802], mem[803], 
        mem[804], mem[805], mem[806], mem[807], mem[808], mem[809], mem[810], 
        mem[811], mem[812], mem[813], mem[814], mem[815], mem[816], mem[817], 
        mem[818], mem[819], mem[820], mem[821], mem[822], mem[823], mem[824], 
        mem[825], mem[826], mem[827], mem[828], mem[829], mem[830], mem[831], 
        mem[832], mem[833], mem[834], mem[835], mem[836], mem[837], mem[838], 
        mem[839]}), .D20({mem[840], mem[841], mem[842], mem[843], mem[844], 
        mem[845], mem[846], mem[847], mem[848], mem[849], mem[850], mem[851], 
        mem[852], mem[853], mem[854], mem[855], mem[856], mem[857], mem[858], 
        mem[859], mem[860], mem[861], mem[862], mem[863], mem[864], mem[865], 
        mem[866], mem[867], mem[868], mem[869], mem[870], mem[871], mem[872], 
        mem[873], mem[874], mem[875], mem[876], mem[877], mem[878], mem[879], 
        mem[880], mem[881]}), .D21({mem[882], mem[883], mem[884], mem[885], 
        mem[886], mem[887], mem[888], mem[889], mem[890], mem[891], mem[892], 
        mem[893], mem[894], mem[895], mem[896], mem[897], mem[898], mem[899], 
        mem[900], mem[901], mem[902], mem[903], mem[904], mem[905], mem[906], 
        mem[907], mem[908], mem[909], mem[910], mem[911], mem[912], mem[913], 
        mem[914], mem[915], mem[916], mem[917], mem[918], mem[919], mem[920], 
        mem[921], mem[922], mem[923]}), .D22({mem[924], mem[925], mem[926], 
        mem[927], mem[928], mem[929], mem[930], mem[931], mem[932], mem[933], 
        mem[934], mem[935], mem[936], mem[937], mem[938], mem[939], mem[940], 
        mem[941], mem[942], mem[943], mem[944], mem[945], mem[946], mem[947], 
        mem[948], mem[949], mem[950], mem[951], mem[952], mem[953], mem[954], 
        mem[955], mem[956], mem[957], mem[958], mem[959], mem[960], mem[961], 
        mem[962], mem[963], mem[964], mem[965]}), .D23({mem[966], mem[967], 
        mem[968], mem[969], mem[970], mem[971], mem[972], mem[973], mem[974], 
        mem[975], mem[976], mem[977], mem[978], mem[979], mem[980], mem[981], 
        mem[982], mem[983], mem[984], mem[985], mem[986], mem[987], mem[988], 
        mem[989], mem[990], mem[991], mem[992], mem[993], mem[994], mem[995], 
        mem[996], mem[997], mem[998], mem[999], mem[1000], mem[1001], 
        mem[1002], mem[1003], mem[1004], mem[1005], mem[1006], mem[1007]}), 
        .D24({mem[1008], mem[1009], mem[1010], mem[1011], mem[1012], mem[1013], 
        mem[1014], mem[1015], mem[1016], mem[1017], mem[1018], mem[1019], 
        mem[1020], mem[1021], mem[1022], mem[1023], mem[1024], mem[1025], 
        mem[1026], mem[1027], mem[1028], mem[1029], mem[1030], mem[1031], 
        mem[1032], mem[1033], mem[1034], mem[1035], mem[1036], mem[1037], 
        mem[1038], mem[1039], mem[1040], mem[1041], mem[1042], mem[1043], 
        mem[1044], mem[1045], mem[1046], mem[1047], mem[1048], mem[1049]}), 
        .D25({mem[1050], mem[1051], mem[1052], mem[1053], mem[1054], mem[1055], 
        mem[1056], mem[1057], mem[1058], mem[1059], mem[1060], mem[1061], 
        mem[1062], mem[1063], mem[1064], mem[1065], mem[1066], mem[1067], 
        mem[1068], mem[1069], mem[1070], mem[1071], mem[1072], mem[1073], 
        mem[1074], mem[1075], mem[1076], mem[1077], mem[1078], mem[1079], 
        mem[1080], mem[1081], mem[1082], mem[1083], mem[1084], mem[1085], 
        mem[1086], mem[1087], mem[1088], mem[1089], mem[1090], mem[1091]}), 
        .D26({mem[1092], mem[1093], mem[1094], mem[1095], mem[1096], mem[1097], 
        mem[1098], mem[1099], mem[1100], mem[1101], mem[1102], mem[1103], 
        mem[1104], mem[1105], mem[1106], mem[1107], mem[1108], mem[1109], 
        mem[1110], mem[1111], mem[1112], mem[1113], mem[1114], mem[1115], 
        mem[1116], mem[1117], mem[1118], mem[1119], mem[1120], mem[1121], 
        mem[1122], mem[1123], mem[1124], mem[1125], mem[1126], mem[1127], 
        mem[1128], mem[1129], mem[1130], mem[1131], mem[1132], mem[1133]}), 
        .D27({mem[1134], mem[1135], mem[1136], mem[1137], mem[1138], mem[1139], 
        mem[1140], mem[1141], mem[1142], mem[1143], mem[1144], mem[1145], 
        mem[1146], mem[1147], mem[1148], mem[1149], mem[1150], mem[1151], 
        mem[1152], mem[1153], mem[1154], mem[1155], mem[1156], mem[1157], 
        mem[1158], mem[1159], mem[1160], mem[1161], mem[1162], mem[1163], 
        mem[1164], mem[1165], mem[1166], mem[1167], mem[1168], mem[1169], 
        mem[1170], mem[1171], mem[1172], mem[1173], mem[1174], mem[1175]}), 
        .D28({mem[1176], mem[1177], mem[1178], mem[1179], mem[1180], mem[1181], 
        mem[1182], mem[1183], mem[1184], mem[1185], mem[1186], mem[1187], 
        mem[1188], mem[1189], mem[1190], mem[1191], mem[1192], mem[1193], 
        mem[1194], mem[1195], mem[1196], mem[1197], mem[1198], mem[1199], 
        mem[1200], mem[1201], mem[1202], mem[1203], mem[1204], mem[1205], 
        mem[1206], mem[1207], mem[1208], mem[1209], mem[1210], mem[1211], 
        mem[1212], mem[1213], mem[1214], mem[1215], mem[1216], mem[1217]}), 
        .D29({mem[1218], mem[1219], mem[1220], mem[1221], mem[1222], mem[1223], 
        mem[1224], mem[1225], mem[1226], mem[1227], mem[1228], mem[1229], 
        mem[1230], mem[1231], mem[1232], mem[1233], mem[1234], mem[1235], 
        mem[1236], mem[1237], mem[1238], mem[1239], mem[1240], mem[1241], 
        mem[1242], mem[1243], mem[1244], mem[1245], mem[1246], mem[1247], 
        mem[1248], mem[1249], mem[1250], mem[1251], mem[1252], mem[1253], 
        mem[1254], mem[1255], mem[1256], mem[1257], mem[1258], mem[1259]}), 
        .D30({mem[1260], mem[1261], mem[1262], mem[1263], mem[1264], mem[1265], 
        mem[1266], mem[1267], mem[1268], mem[1269], mem[1270], mem[1271], 
        mem[1272], mem[1273], mem[1274], mem[1275], mem[1276], mem[1277], 
        mem[1278], mem[1279], mem[1280], mem[1281], mem[1282], mem[1283], 
        mem[1284], mem[1285], mem[1286], mem[1287], mem[1288], mem[1289], 
        mem[1290], mem[1291], mem[1292], mem[1293], mem[1294], mem[1295], 
        mem[1296], mem[1297], mem[1298], mem[1299], mem[1300], mem[1301]}), 
        .D31({mem[1302], mem[1303], mem[1304], mem[1305], mem[1306], mem[1307], 
        mem[1308], mem[1309], mem[1310], mem[1311], mem[1312], mem[1313], 
        mem[1314], mem[1315], mem[1316], mem[1317], mem[1318], mem[1319], 
        mem[1320], mem[1321], mem[1322], mem[1323], mem[1324], mem[1325], 
        mem[1326], mem[1327], mem[1328], mem[1329], mem[1330], mem[1331], 
        mem[1332], mem[1333], mem[1334], mem[1335], mem[1336], mem[1337], 
        mem[1338], mem[1339], mem[1340], mem[1341], mem[1342], mem[1343]}), 
        .S0(N18), .S1(N19), .S2(N20), .S3(N21), .S4(N22), .Z({data_out[0], 
        data_out[1], data_out[2], data_out[3], data_out[4], data_out[5], 
        data_out[6], data_out[7], data_out[8], data_out[9], data_out[10], 
        data_out[11], data_out[12], data_out[13], data_out[14], data_out[15], 
        data_out[16], data_out[17], data_out[18], data_out[19], data_out[20], 
        data_out[21], data_out[22], data_out[23], data_out[24], data_out[25], 
        data_out[26], data_out[27], data_out[28], data_out[29], data_out[30], 
        data_out[31], data_out[32], data_out[33], data_out[34], data_out[35], 
        data_out[36], data_out[37], data_out[38], data_out[39], data_out[40], 
        data_out[41]}) );
  GTECH_BUF B_2 ( .A(rd_ptr[0]), .Z(N18) );
  GTECH_BUF B_3 ( .A(rd_ptr[1]), .Z(N19) );
  GTECH_BUF B_4 ( .A(rd_ptr[2]), .Z(N20) );
  GTECH_BUF B_5 ( .A(rd_ptr[3]), .Z(N21) );
  GTECH_BUF B_6 ( .A(rd_ptr[4]), .Z(N22) );
  GTECH_AND2 C11258 ( .A(N228), .B(put), .Z(N23) );
  GTECH_NOT I_18 ( .A(fillcount[5]), .Z(N228) );
  GTECH_AND2 C11261 ( .A(N229), .B(get), .Z(N24) );
  GTECH_AND2 C11262 ( .A(N23), .B(N128), .Z(N229) );
  GTECH_AND2 C11263 ( .A(N128), .B(get), .Z(N25) );
  GTECH_OR2 C11268 ( .A(N24), .B(reset), .Z(N26) );
  GTECH_OR2 C11269 ( .A(N23), .B(N26), .Z(N27) );
  GTECH_OR2 C11270 ( .A(N25), .B(N27), .Z(N28) );
  GTECH_NOT I_19 ( .A(N28), .Z(N29) );
  GTECH_BUF B_7 ( .A(N117), .Z(N30) );
  GTECH_BUF B_8 ( .A(N120), .Z(N41) );
  GTECH_BUF B_9 ( .A(N123), .Z(N53) );
  GTECH_NOT I_20 ( .A(reset), .Z(N116) );
  GTECH_AND2 C11340 ( .A(N24), .B(N116), .Z(N117) );
  GTECH_AND2 C11341 ( .A(N30), .B(N116), .Z(net421) );
  GTECH_NOT I_21 ( .A(N24), .Z(N118) );
  GTECH_AND2 C11343 ( .A(N116), .B(N118), .Z(N119) );
  GTECH_AND2 C11344 ( .A(N23), .B(N119), .Z(N120) );
  GTECH_AND2 C11345 ( .A(N41), .B(N119), .Z(net422) );
  GTECH_NOT I_22 ( .A(N23), .Z(N121) );
  GTECH_AND2 C11347 ( .A(N119), .B(N121), .Z(N122) );
  GTECH_AND2 C11348 ( .A(N25), .B(N122), .Z(N123) );
  GTECH_AND2 C11349 ( .A(N53), .B(N122), .Z(net423) );
endmodule


module ddr3_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, dm, odt, 
        ts_con, cke, resetbar, clk, reset, init, ck );
  output [2:0] ba;
  output [13:0] a;
  output [1:0] dm;
  input clk, reset, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke, resetbar;
  wire   N0, N1, N2, N3, flag, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14,
         N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         net500;
  wire   [18:0] counter;
  tri   ready;
  tri   clk;
  tri   reset;
  tri   ck;

  GTECH_AND2 C22 ( .A(N29), .B(N30), .Z(N31) );
  GTECH_AND2 C43 ( .A(N33), .B(N34), .Z(N50) );
  GTECH_AND2 C44 ( .A(N35), .B(N36), .Z(N51) );
  GTECH_AND2 C45 ( .A(N37), .B(N38), .Z(N52) );
  GTECH_AND2 C46 ( .A(N39), .B(N40), .Z(N53) );
  GTECH_AND2 C47 ( .A(N41), .B(N42), .Z(N54) );
  GTECH_AND2 C48 ( .A(N43), .B(N44), .Z(N55) );
  GTECH_AND2 C49 ( .A(N45), .B(N46), .Z(N56) );
  GTECH_AND2 C50 ( .A(N47), .B(N48), .Z(N57) );
  GTECH_AND2 C51 ( .A(N50), .B(N51), .Z(N58) );
  GTECH_AND2 C52 ( .A(N52), .B(N53), .Z(N59) );
  GTECH_AND2 C53 ( .A(N54), .B(N55), .Z(N60) );
  GTECH_AND2 C54 ( .A(N56), .B(N57), .Z(N61) );
  GTECH_AND2 C55 ( .A(N58), .B(N59), .Z(N62) );
  GTECH_AND2 C56 ( .A(N60), .B(N61), .Z(N63) );
  GTECH_AND2 C57 ( .A(N62), .B(N63), .Z(N64) );
  GTECH_AND2 C58 ( .A(N64), .B(N49), .Z(N65) );
  GTECH_OR2 C66 ( .A(counter[17]), .B(counter[16]), .Z(N66) );
  GTECH_OR2 C67 ( .A(N35), .B(N36), .Z(N67) );
  GTECH_OR2 C68 ( .A(N37), .B(N38), .Z(N68) );
  GTECH_OR2 C69 ( .A(counter[11]), .B(N40), .Z(N69) );
  GTECH_OR2 C70 ( .A(counter[9]), .B(counter[7]), .Z(N70) );
  GTECH_OR2 C71 ( .A(counter[6]), .B(N44), .Z(N71) );
  GTECH_OR2 C72 ( .A(counter[4]), .B(counter[3]), .Z(N72) );
  GTECH_OR2 C73 ( .A(N47), .B(counter[1]), .Z(N73) );
  GTECH_OR2 C74 ( .A(N66), .B(N67), .Z(N74) );
  GTECH_OR2 C75 ( .A(N68), .B(N69), .Z(N75) );
  GTECH_OR2 C76 ( .A(N70), .B(N71), .Z(N76) );
  GTECH_OR2 C77 ( .A(N72), .B(N73), .Z(N77) );
  GTECH_OR2 C78 ( .A(N74), .B(N75), .Z(N78) );
  GTECH_OR2 C79 ( .A(N76), .B(N77), .Z(N79) );
  GTECH_OR2 C80 ( .A(N78), .B(N79), .Z(N80) );
  GTECH_OR2 C81 ( .A(N80), .B(counter[0]), .Z(N81) );
  GTECH_OR2 C90 ( .A(counter[17]), .B(counter[16]), .Z(N83) );
  GTECH_OR2 C91 ( .A(N35), .B(N36), .Z(N84) );
  GTECH_OR2 C92 ( .A(N37), .B(N38), .Z(N85) );
  GTECH_OR2 C93 ( .A(counter[11]), .B(N40), .Z(N86) );
  GTECH_OR2 C94 ( .A(counter[9]), .B(counter[7]), .Z(N87) );
  GTECH_OR2 C95 ( .A(counter[6]), .B(N44), .Z(N88) );
  GTECH_OR2 C96 ( .A(counter[4]), .B(N46), .Z(N89) );
  GTECH_OR2 C97 ( .A(counter[2]), .B(counter[1]), .Z(N90) );
  GTECH_OR2 C98 ( .A(N83), .B(N84), .Z(N91) );
  GTECH_OR2 C99 ( .A(N85), .B(N86), .Z(N92) );
  GTECH_OR2 C100 ( .A(N87), .B(N88), .Z(N93) );
  GTECH_OR2 C101 ( .A(N89), .B(N90), .Z(N94) );
  GTECH_OR2 C102 ( .A(N91), .B(N92), .Z(N95) );
  GTECH_OR2 C103 ( .A(N93), .B(N94), .Z(N96) );
  GTECH_OR2 C104 ( .A(N95), .B(N96), .Z(N97) );
  GTECH_OR2 C105 ( .A(N97), .B(counter[0]), .Z(N98) );
  GTECH_OR2 C115 ( .A(N33), .B(N34), .Z(N100) );
  GTECH_OR2 C116 ( .A(counter[15]), .B(N36), .Z(N101) );
  GTECH_OR2 C117 ( .A(counter[13]), .B(N38), .Z(N102) );
  GTECH_OR2 C118 ( .A(counter[11]), .B(N40), .Z(N103) );
  GTECH_OR2 C119 ( .A(N41), .B(N42), .Z(N104) );
  GTECH_OR2 C120 ( .A(counter[6]), .B(counter[5]), .Z(N105) );
  GTECH_OR2 C121 ( .A(counter[4]), .B(counter[3]), .Z(N106) );
  GTECH_OR2 C122 ( .A(counter[2]), .B(N48), .Z(N107) );
  GTECH_OR2 C123 ( .A(N100), .B(N101), .Z(N108) );
  GTECH_OR2 C124 ( .A(N102), .B(N103), .Z(N109) );
  GTECH_OR2 C125 ( .A(N104), .B(N105), .Z(N110) );
  GTECH_OR2 C126 ( .A(N106), .B(N107), .Z(N111) );
  GTECH_OR2 C127 ( .A(N108), .B(N109), .Z(N112) );
  GTECH_OR2 C128 ( .A(N110), .B(N111), .Z(N113) );
  GTECH_OR2 C129 ( .A(N112), .B(N113), .Z(N114) );
  GTECH_OR2 C130 ( .A(N114), .B(counter[0]), .Z(N115) );
  GTECH_OR2 C141 ( .A(N33), .B(N34), .Z(N117) );
  GTECH_OR2 C142 ( .A(counter[15]), .B(N36), .Z(N118) );
  GTECH_OR2 C143 ( .A(counter[13]), .B(N38), .Z(N119) );
  GTECH_OR2 C144 ( .A(counter[11]), .B(N40), .Z(N120) );
  GTECH_OR2 C145 ( .A(N41), .B(N42), .Z(N121) );
  GTECH_OR2 C146 ( .A(counter[6]), .B(N44), .Z(N122) );
  GTECH_OR2 C147 ( .A(counter[4]), .B(N46), .Z(N123) );
  GTECH_OR2 C148 ( .A(counter[2]), .B(counter[1]), .Z(N124) );
  GTECH_OR2 C149 ( .A(N117), .B(N118), .Z(N125) );
  GTECH_OR2 C150 ( .A(N119), .B(N120), .Z(N126) );
  GTECH_OR2 C151 ( .A(N121), .B(N122), .Z(N127) );
  GTECH_OR2 C152 ( .A(N123), .B(N124), .Z(N128) );
  GTECH_OR2 C153 ( .A(N125), .B(N126), .Z(N129) );
  GTECH_OR2 C154 ( .A(N127), .B(N128), .Z(N130) );
  GTECH_OR2 C155 ( .A(N129), .B(N130), .Z(N131) );
  GTECH_OR2 C156 ( .A(N131), .B(counter[0]), .Z(N132) );
  GTECH_OR2 C168 ( .A(N33), .B(N34), .Z(N134) );
  GTECH_OR2 C169 ( .A(counter[15]), .B(N36), .Z(N135) );
  GTECH_OR2 C170 ( .A(counter[13]), .B(N38), .Z(N136) );
  GTECH_OR2 C171 ( .A(counter[11]), .B(N40), .Z(N137) );
  GTECH_OR2 C172 ( .A(N41), .B(N42), .Z(N138) );
  GTECH_OR2 C173 ( .A(counter[6]), .B(N44), .Z(N139) );
  GTECH_OR2 C174 ( .A(counter[4]), .B(N46), .Z(N140) );
  GTECH_OR2 C175 ( .A(counter[2]), .B(counter[1]), .Z(N141) );
  GTECH_OR2 C176 ( .A(N134), .B(N135), .Z(N142) );
  GTECH_OR2 C177 ( .A(N136), .B(N137), .Z(N143) );
  GTECH_OR2 C178 ( .A(N138), .B(N139), .Z(N144) );
  GTECH_OR2 C179 ( .A(N140), .B(N141), .Z(N145) );
  GTECH_OR2 C180 ( .A(N142), .B(N143), .Z(N146) );
  GTECH_OR2 C181 ( .A(N144), .B(N145), .Z(N147) );
  GTECH_OR2 C182 ( .A(N146), .B(N147), .Z(N148) );
  GTECH_OR2 C183 ( .A(N148), .B(N49), .Z(N149) );
  GTECH_OR2 C195 ( .A(N33), .B(N34), .Z(N151) );
  GTECH_OR2 C196 ( .A(counter[15]), .B(N36), .Z(N152) );
  GTECH_OR2 C197 ( .A(counter[13]), .B(N38), .Z(N153) );
  GTECH_OR2 C198 ( .A(counter[11]), .B(N40), .Z(N154) );
  GTECH_OR2 C199 ( .A(N41), .B(N42), .Z(N155) );
  GTECH_OR2 C200 ( .A(counter[6]), .B(N44), .Z(N156) );
  GTECH_OR2 C201 ( .A(counter[4]), .B(N46), .Z(N157) );
  GTECH_OR2 C202 ( .A(N47), .B(counter[1]), .Z(N158) );
  GTECH_OR2 C203 ( .A(N151), .B(N152), .Z(N159) );
  GTECH_OR2 C204 ( .A(N153), .B(N154), .Z(N160) );
  GTECH_OR2 C205 ( .A(N155), .B(N156), .Z(N161) );
  GTECH_OR2 C206 ( .A(N157), .B(N158), .Z(N162) );
  GTECH_OR2 C207 ( .A(N159), .B(N160), .Z(N163) );
  GTECH_OR2 C208 ( .A(N161), .B(N162), .Z(N164) );
  GTECH_OR2 C209 ( .A(N163), .B(N164), .Z(N165) );
  GTECH_OR2 C210 ( .A(N165), .B(counter[0]), .Z(N166) );
  GTECH_OR2 C223 ( .A(N33), .B(N34), .Z(N168) );
  GTECH_OR2 C224 ( .A(counter[15]), .B(N36), .Z(N169) );
  GTECH_OR2 C225 ( .A(counter[13]), .B(N38), .Z(N170) );
  GTECH_OR2 C226 ( .A(counter[11]), .B(N40), .Z(N171) );
  GTECH_OR2 C227 ( .A(N41), .B(N42), .Z(N172) );
  GTECH_OR2 C228 ( .A(counter[6]), .B(N44), .Z(N173) );
  GTECH_OR2 C229 ( .A(counter[4]), .B(N46), .Z(N174) );
  GTECH_OR2 C230 ( .A(N47), .B(counter[1]), .Z(N175) );
  GTECH_OR2 C231 ( .A(N168), .B(N169), .Z(N176) );
  GTECH_OR2 C232 ( .A(N170), .B(N171), .Z(N177) );
  GTECH_OR2 C233 ( .A(N172), .B(N173), .Z(N178) );
  GTECH_OR2 C234 ( .A(N174), .B(N175), .Z(N179) );
  GTECH_OR2 C235 ( .A(N176), .B(N177), .Z(N180) );
  GTECH_OR2 C236 ( .A(N178), .B(N179), .Z(N181) );
  GTECH_OR2 C237 ( .A(N180), .B(N181), .Z(N182) );
  GTECH_OR2 C238 ( .A(N182), .B(N49), .Z(N183) );
  GTECH_OR2 C249 ( .A(N33), .B(N34), .Z(N185) );
  GTECH_OR2 C250 ( .A(counter[15]), .B(N36), .Z(N186) );
  GTECH_OR2 C251 ( .A(counter[13]), .B(N38), .Z(N187) );
  GTECH_OR2 C252 ( .A(counter[11]), .B(N40), .Z(N188) );
  GTECH_OR2 C253 ( .A(N41), .B(N42), .Z(N189) );
  GTECH_OR2 C254 ( .A(counter[6]), .B(N44), .Z(N190) );
  GTECH_OR2 C255 ( .A(N45), .B(counter[3]), .Z(N191) );
  GTECH_OR2 C256 ( .A(counter[2]), .B(counter[1]), .Z(N192) );
  GTECH_OR2 C257 ( .A(N185), .B(N186), .Z(N193) );
  GTECH_OR2 C258 ( .A(N187), .B(N188), .Z(N194) );
  GTECH_OR2 C259 ( .A(N189), .B(N190), .Z(N195) );
  GTECH_OR2 C260 ( .A(N191), .B(N192), .Z(N196) );
  GTECH_OR2 C261 ( .A(N193), .B(N194), .Z(N197) );
  GTECH_OR2 C262 ( .A(N195), .B(N196), .Z(N198) );
  GTECH_OR2 C263 ( .A(N197), .B(N198), .Z(N199) );
  GTECH_OR2 C264 ( .A(N199), .B(counter[0]), .Z(N200) );
  GTECH_OR2 C276 ( .A(N33), .B(N34), .Z(N202) );
  GTECH_OR2 C277 ( .A(counter[15]), .B(N36), .Z(N203) );
  GTECH_OR2 C278 ( .A(counter[13]), .B(N38), .Z(N204) );
  GTECH_OR2 C279 ( .A(counter[11]), .B(N40), .Z(N205) );
  GTECH_OR2 C280 ( .A(N41), .B(N42), .Z(N206) );
  GTECH_OR2 C281 ( .A(counter[6]), .B(N44), .Z(N207) );
  GTECH_OR2 C282 ( .A(N45), .B(counter[3]), .Z(N208) );
  GTECH_OR2 C283 ( .A(counter[2]), .B(counter[1]), .Z(N209) );
  GTECH_OR2 C284 ( .A(N202), .B(N203), .Z(N210) );
  GTECH_OR2 C285 ( .A(N204), .B(N205), .Z(N211) );
  GTECH_OR2 C286 ( .A(N206), .B(N207), .Z(N212) );
  GTECH_OR2 C287 ( .A(N208), .B(N209), .Z(N213) );
  GTECH_OR2 C288 ( .A(N210), .B(N211), .Z(N214) );
  GTECH_OR2 C289 ( .A(N212), .B(N213), .Z(N215) );
  GTECH_OR2 C290 ( .A(N214), .B(N215), .Z(N216) );
  GTECH_OR2 C291 ( .A(N216), .B(N49), .Z(N217) );
  GTECH_OR2 C303 ( .A(N33), .B(N34), .Z(N219) );
  GTECH_OR2 C304 ( .A(counter[15]), .B(N36), .Z(N220) );
  GTECH_OR2 C305 ( .A(counter[13]), .B(N38), .Z(N221) );
  GTECH_OR2 C306 ( .A(counter[11]), .B(N40), .Z(N222) );
  GTECH_OR2 C307 ( .A(N41), .B(N42), .Z(N223) );
  GTECH_OR2 C308 ( .A(counter[6]), .B(N44), .Z(N224) );
  GTECH_OR2 C309 ( .A(N45), .B(counter[3]), .Z(N225) );
  GTECH_OR2 C310 ( .A(N47), .B(counter[1]), .Z(N226) );
  GTECH_OR2 C311 ( .A(N219), .B(N220), .Z(N227) );
  GTECH_OR2 C312 ( .A(N221), .B(N222), .Z(N228) );
  GTECH_OR2 C313 ( .A(N223), .B(N224), .Z(N229) );
  GTECH_OR2 C314 ( .A(N225), .B(N226), .Z(N230) );
  GTECH_OR2 C315 ( .A(N227), .B(N228), .Z(N231) );
  GTECH_OR2 C316 ( .A(N229), .B(N230), .Z(N232) );
  GTECH_OR2 C317 ( .A(N231), .B(N232), .Z(N233) );
  GTECH_OR2 C318 ( .A(N233), .B(counter[0]), .Z(N234) );
  GTECH_OR2 C331 ( .A(N33), .B(N34), .Z(N236) );
  GTECH_OR2 C332 ( .A(counter[15]), .B(N36), .Z(N237) );
  GTECH_OR2 C333 ( .A(counter[13]), .B(N38), .Z(N238) );
  GTECH_OR2 C334 ( .A(counter[11]), .B(N40), .Z(N239) );
  GTECH_OR2 C335 ( .A(N41), .B(N42), .Z(N240) );
  GTECH_OR2 C336 ( .A(counter[6]), .B(N44), .Z(N241) );
  GTECH_OR2 C337 ( .A(N45), .B(counter[3]), .Z(N242) );
  GTECH_OR2 C338 ( .A(N47), .B(counter[1]), .Z(N243) );
  GTECH_OR2 C339 ( .A(N236), .B(N237), .Z(N244) );
  GTECH_OR2 C340 ( .A(N238), .B(N239), .Z(N245) );
  GTECH_OR2 C341 ( .A(N240), .B(N241), .Z(N246) );
  GTECH_OR2 C342 ( .A(N242), .B(N243), .Z(N247) );
  GTECH_OR2 C343 ( .A(N244), .B(N245), .Z(N248) );
  GTECH_OR2 C344 ( .A(N246), .B(N247), .Z(N249) );
  GTECH_OR2 C345 ( .A(N248), .B(N249), .Z(N250) );
  GTECH_OR2 C346 ( .A(N250), .B(N49), .Z(N251) );
  GTECH_OR2 C356 ( .A(N33), .B(N34), .Z(N253) );
  GTECH_OR2 C357 ( .A(counter[15]), .B(N36), .Z(N254) );
  GTECH_OR2 C358 ( .A(counter[13]), .B(N38), .Z(N255) );
  GTECH_OR2 C359 ( .A(counter[11]), .B(N40), .Z(N256) );
  GTECH_OR2 C360 ( .A(N41), .B(N42), .Z(N257) );
  GTECH_OR2 C361 ( .A(N43), .B(counter[5]), .Z(N258) );
  GTECH_OR2 C362 ( .A(counter[4]), .B(counter[3]), .Z(N259) );
  GTECH_OR2 C363 ( .A(counter[2]), .B(counter[1]), .Z(N260) );
  GTECH_OR2 C364 ( .A(N253), .B(N254), .Z(N261) );
  GTECH_OR2 C365 ( .A(N255), .B(N256), .Z(N262) );
  GTECH_OR2 C366 ( .A(N257), .B(N258), .Z(N263) );
  GTECH_OR2 C367 ( .A(N259), .B(N260), .Z(N264) );
  GTECH_OR2 C368 ( .A(N261), .B(N262), .Z(N265) );
  GTECH_OR2 C369 ( .A(N263), .B(N264), .Z(N266) );
  GTECH_OR2 C370 ( .A(N265), .B(N266), .Z(N267) );
  GTECH_OR2 C371 ( .A(N267), .B(counter[0]), .Z(N268) );
  GTECH_OR2 C382 ( .A(N33), .B(N34), .Z(N270) );
  GTECH_OR2 C383 ( .A(counter[15]), .B(N36), .Z(N271) );
  GTECH_OR2 C384 ( .A(counter[13]), .B(N38), .Z(N272) );
  GTECH_OR2 C385 ( .A(counter[11]), .B(N40), .Z(N273) );
  GTECH_OR2 C386 ( .A(N41), .B(N42), .Z(N274) );
  GTECH_OR2 C387 ( .A(N43), .B(counter[5]), .Z(N275) );
  GTECH_OR2 C388 ( .A(counter[4]), .B(counter[3]), .Z(N276) );
  GTECH_OR2 C389 ( .A(counter[2]), .B(counter[1]), .Z(N277) );
  GTECH_OR2 C390 ( .A(N270), .B(N271), .Z(N278) );
  GTECH_OR2 C391 ( .A(N272), .B(N273), .Z(N279) );
  GTECH_OR2 C392 ( .A(N274), .B(N275), .Z(N280) );
  GTECH_OR2 C393 ( .A(N276), .B(N277), .Z(N281) );
  GTECH_OR2 C394 ( .A(N278), .B(N279), .Z(N282) );
  GTECH_OR2 C395 ( .A(N280), .B(N281), .Z(N283) );
  GTECH_OR2 C396 ( .A(N282), .B(N283), .Z(N284) );
  GTECH_OR2 C397 ( .A(N284), .B(N49), .Z(N285) );
  GTECH_OR2 C407 ( .A(N33), .B(N34), .Z(N287) );
  GTECH_OR2 C408 ( .A(counter[15]), .B(N36), .Z(N288) );
  GTECH_OR2 C409 ( .A(counter[13]), .B(N38), .Z(N289) );
  GTECH_OR2 C410 ( .A(N39), .B(counter[10]), .Z(N290) );
  GTECH_OR2 C411 ( .A(counter[9]), .B(N42), .Z(N291) );
  GTECH_OR2 C412 ( .A(N43), .B(counter[5]), .Z(N292) );
  GTECH_OR2 C413 ( .A(counter[4]), .B(counter[3]), .Z(N293) );
  GTECH_OR2 C414 ( .A(counter[2]), .B(counter[1]), .Z(N294) );
  GTECH_OR2 C415 ( .A(N287), .B(N288), .Z(N295) );
  GTECH_OR2 C416 ( .A(N289), .B(N290), .Z(N296) );
  GTECH_OR2 C417 ( .A(N291), .B(N292), .Z(N297) );
  GTECH_OR2 C418 ( .A(N293), .B(N294), .Z(N298) );
  GTECH_OR2 C419 ( .A(N295), .B(N296), .Z(N299) );
  GTECH_OR2 C420 ( .A(N297), .B(N298), .Z(N300) );
  GTECH_OR2 C421 ( .A(N299), .B(N300), .Z(N301) );
  GTECH_OR2 C422 ( .A(N301), .B(N49), .Z(N302) );
  \**SEQGEN**  rasbar_reg ( .clear(1'b0), .preset(1'b0), .next_state(N348), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(rasbar), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N346) );
  \**SEQGEN**  webar_reg ( .clear(1'b0), .preset(1'b0), .next_state(N347), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(webar), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N346) );
  \**SEQGEN**  casbar_reg ( .clear(1'b0), .preset(1'b0), .next_state(N348), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(casbar), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N346) );
  \**SEQGEN**  ready_reg ( .clear(1'b0), .preset(1'b0), .next_state(N350), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ready), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N349) );
  \**SEQGEN**  counter_reg_18_ ( .clear(1'b0), .preset(1'b0), .next_state(N371), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_17_ ( .clear(1'b0), .preset(1'b0), .next_state(N370), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_16_ ( .clear(1'b0), .preset(1'b0), .next_state(N369), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_15_ ( .clear(1'b0), .preset(1'b0), .next_state(N368), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_14_ ( .clear(1'b0), .preset(1'b0), .next_state(N367), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(N366), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(N365), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(N364), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(N363), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(N362), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(N361), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(N360), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(N359), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N358), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N357), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N356), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N355), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N354), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  counter_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N353), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(counter[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N372) );
  \**SEQGEN**  resetbar_reg ( .clear(1'b0), .preset(1'b0), .next_state(N352), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(resetbar), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N351) );
  \**SEQGEN**  flag_reg ( .clear(1'b0), .preset(1'b0), .next_state(N372), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(flag), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N336) );
  \**SEQGEN**  cke_reg ( .clear(1'b0), .preset(1'b0), .next_state(N338), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(cke), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N337) );
  \**SEQGEN**  odt_reg ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(odt), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(reset) );
  \**SEQGEN**  a_reg_13_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_12_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_11_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(N342), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(N340), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(N340), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N341), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N340), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  a_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(a[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N339) );
  \**SEQGEN**  ba_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ba[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N343) );
  \**SEQGEN**  ba_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N345), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ba[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N343) );
  \**SEQGEN**  ba_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N344), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ba[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N343) );
  \**SEQGEN**  ts_con_reg ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ts_con), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(reset) );
  \**SEQGEN**  csbar_reg ( .clear(1'b0), .preset(1'b0), .next_state(N347), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(csbar), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N346) );
  GTECH_NOT I_0 ( .A(flag), .Z(N377) );
  GTECH_OR2 C704 ( .A(N374), .B(N350), .Z(N372) );
  GTECH_OR2 C707 ( .A(N167), .B(N201), .Z(N324) );
  GTECH_OR2 C709 ( .A(N133), .B(N167), .Z(N325) );
  GTECH_OR2 C710 ( .A(N201), .B(N235), .Z(N327) );
  GTECH_OR4 C721 ( .A(N133), .B(N167), .C(N201), .D(N235), .Z(N323) );
  GTECH_OR5 C723 ( .A(N82), .B(N116), .C(N150), .D(N184), .E(N218), .Z(N378)
         );
  GTECH_OR2 C724 ( .A(N252), .B(N286), .Z(N379) );
  GTECH_OR2 C725 ( .A(N378), .B(N379), .Z(N320) );
  GTECH_OR5 C726 ( .A(N133), .B(N167), .C(N201), .D(N235), .E(N269), .Z(N326)
         );
  GTECH_OR3 C734 ( .A(N252), .B(N269), .C(N286), .Z(N380) );
  GTECH_OR2 C735 ( .A(N378), .B(N380), .Z(N321) );
  ADD_UNS_OP add_90 ( .A(counter), .B(1'b1), .Z({N28, N27, N26, N25, N24, N23, 
        N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10}) );
  GTECH_OR2 C762 ( .A(N65), .B(N99), .Z(N318) );
  GTECH_OR5 C763 ( .A(N82), .B(N116), .C(N133), .D(N150), .E(N167), .Z(N381)
         );
  GTECH_OR5 C764 ( .A(N184), .B(N201), .C(N218), .D(N235), .E(N252), .Z(N382)
         );
  GTECH_OR2 C771 ( .A(N269), .B(N286), .Z(N383) );
  GTECH_OR3 C772 ( .A(N381), .B(N382), .C(N383), .Z(N319) );
  GTECH_OR2 C796 ( .A(N82), .B(N116), .Z(N322) );
  GTECH_OR2 C896 ( .A(N374), .B(N8), .Z(N384) );
  GTECH_OR2 C944 ( .A(reset), .B(N374), .Z(N385) );
  GTECH_NOT I_1 ( .A(N317), .Z(N328) );
  SELECT_OP C949 ( .DATA1(N303), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N329) );
  GTECH_BUF B_0 ( .A(N31), .Z(N0) );
  SELECT_OP C950 ( .DATA1(N328), .DATA2(1'b1), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N330) );
  SELECT_OP C951 ( .DATA1(N318), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N331) );
  SELECT_OP C952 ( .DATA1(N319), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N332) );
  SELECT_OP C953 ( .DATA1(N322), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N333) );
  SELECT_OP C954 ( .DATA1(N323), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N334) );
  SELECT_OP C955 ( .DATA1(N326), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N32), 
        .Z(N335) );
  SELECT_OP C956 ( .DATA1(1'b1), .DATA2(N330), .DATA3(1'b0), .CONTROL1(N1), 
        .CONTROL2(N350), .CONTROL3(N8), .Z(N336) );
  GTECH_BUF B_1 ( .A(N385), .Z(N1) );
  SELECT_OP C957 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N333), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N337) );
  GTECH_BUF B_2 ( .A(reset), .Z(N2) );
  GTECH_BUF B_3 ( .A(N384), .Z(N3) );
  SELECT_OP C958 ( .DATA1(1'b0), .DATA2(N116), .CONTROL1(N2), .CONTROL2(N350), 
        .Z(N338) );
  SELECT_OP C959 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N335), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N339) );
  SELECT_OP C960 ( .DATA1({1'b0, 1'b0, 1'b0}), .DATA2({N269, N327, N235}), 
        .CONTROL1(N2), .CONTROL2(N350), .Z({N342, N341, N340}) );
  SELECT_OP C961 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N334), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N343) );
  SELECT_OP C962 ( .DATA1({1'b0, 1'b0}), .DATA2({N325, N324}), .CONTROL1(N2), 
        .CONTROL2(N350), .Z({N345, N344}) );
  SELECT_OP C963 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N332), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N346) );
  SELECT_OP C964 ( .DATA1(1'b1), .DATA2(N320), .CONTROL1(N2), .CONTROL2(N350), 
        .Z(N347) );
  SELECT_OP C965 ( .DATA1(1'b1), .DATA2(N321), .CONTROL1(N2), .CONTROL2(N350), 
        .Z(N348) );
  SELECT_OP C966 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N329), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N349) );
  SELECT_OP C967 ( .DATA1(1'b1), .DATA2(1'b0), .DATA3(N331), .CONTROL1(N2), 
        .CONTROL2(N3), .CONTROL3(N350), .Z(N351) );
  SELECT_OP C968 ( .DATA1(1'b0), .DATA2(N99), .CONTROL1(N2), .CONTROL2(N350), 
        .Z(N352) );
  SELECT_OP C969 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2({N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10}), .CONTROL1(N374), .CONTROL2(N350), 
        .Z({N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353}) );
  GTECH_AND2 C972 ( .A(N377), .B(init), .Z(N4) );
  GTECH_AND2 C973 ( .A(flag), .B(ck), .Z(N5) );
  GTECH_OR2 C977 ( .A(N4), .B(reset), .Z(N6) );
  GTECH_OR2 C978 ( .A(N5), .B(N6), .Z(N7) );
  GTECH_NOT I_2 ( .A(N7), .Z(N8) );
  GTECH_BUF B_4 ( .A(N350), .Z(N9) );
  GTECH_NOT I_3 ( .A(counter[18]), .Z(N29) );
  GTECH_NOT I_4 ( .A(counter[8]), .Z(N30) );
  GTECH_NOT I_5 ( .A(N31), .Z(N32) );
  GTECH_NOT I_6 ( .A(counter[17]), .Z(N33) );
  GTECH_NOT I_7 ( .A(counter[16]), .Z(N34) );
  GTECH_NOT I_8 ( .A(counter[15]), .Z(N35) );
  GTECH_NOT I_9 ( .A(counter[14]), .Z(N36) );
  GTECH_NOT I_10 ( .A(counter[13]), .Z(N37) );
  GTECH_NOT I_11 ( .A(counter[12]), .Z(N38) );
  GTECH_NOT I_12 ( .A(counter[11]), .Z(N39) );
  GTECH_NOT I_13 ( .A(counter[10]), .Z(N40) );
  GTECH_NOT I_14 ( .A(counter[9]), .Z(N41) );
  GTECH_NOT I_15 ( .A(counter[7]), .Z(N42) );
  GTECH_NOT I_16 ( .A(counter[6]), .Z(N43) );
  GTECH_NOT I_17 ( .A(counter[5]), .Z(N44) );
  GTECH_NOT I_18 ( .A(counter[4]), .Z(N45) );
  GTECH_NOT I_19 ( .A(counter[3]), .Z(N46) );
  GTECH_NOT I_20 ( .A(counter[2]), .Z(N47) );
  GTECH_NOT I_21 ( .A(counter[1]), .Z(N48) );
  GTECH_NOT I_22 ( .A(counter[0]), .Z(N49) );
  GTECH_NOT I_23 ( .A(N81), .Z(N82) );
  GTECH_NOT I_24 ( .A(N98), .Z(N99) );
  GTECH_NOT I_25 ( .A(N115), .Z(N116) );
  GTECH_NOT I_26 ( .A(N132), .Z(N133) );
  GTECH_NOT I_27 ( .A(N149), .Z(N150) );
  GTECH_NOT I_28 ( .A(N166), .Z(N167) );
  GTECH_NOT I_29 ( .A(N183), .Z(N184) );
  GTECH_NOT I_30 ( .A(N200), .Z(N201) );
  GTECH_NOT I_31 ( .A(N217), .Z(N218) );
  GTECH_NOT I_32 ( .A(N234), .Z(N235) );
  GTECH_NOT I_33 ( .A(N251), .Z(N252) );
  GTECH_NOT I_34 ( .A(N268), .Z(N269) );
  GTECH_NOT I_35 ( .A(N285), .Z(N286) );
  GTECH_NOT I_36 ( .A(N302), .Z(N303) );
  GTECH_OR2 C1158 ( .A(N82), .B(N65), .Z(N304) );
  GTECH_OR2 C1159 ( .A(N99), .B(N304), .Z(N305) );
  GTECH_OR2 C1160 ( .A(N116), .B(N305), .Z(N306) );
  GTECH_OR2 C1161 ( .A(N133), .B(N306), .Z(N307) );
  GTECH_OR2 C1162 ( .A(N150), .B(N307), .Z(N308) );
  GTECH_OR2 C1163 ( .A(N167), .B(N308), .Z(N309) );
  GTECH_OR2 C1164 ( .A(N184), .B(N309), .Z(N310) );
  GTECH_OR2 C1165 ( .A(N201), .B(N310), .Z(N311) );
  GTECH_OR2 C1166 ( .A(N218), .B(N311), .Z(N312) );
  GTECH_OR2 C1167 ( .A(N235), .B(N312), .Z(N313) );
  GTECH_OR2 C1168 ( .A(N252), .B(N313), .Z(N314) );
  GTECH_OR2 C1169 ( .A(N269), .B(N314), .Z(N315) );
  GTECH_OR2 C1170 ( .A(N286), .B(N315), .Z(N316) );
  GTECH_OR2 C1171 ( .A(N303), .B(N316), .Z(N317) );
  GTECH_NOT I_37 ( .A(reset), .Z(N373) );
  GTECH_AND2 C1174 ( .A(N4), .B(N373), .Z(N374) );
  GTECH_NOT I_38 ( .A(N4), .Z(N375) );
  GTECH_AND2 C1176 ( .A(N373), .B(N375), .Z(N376) );
  GTECH_AND2 C1177 ( .A(N5), .B(N376), .Z(N350) );
  GTECH_AND2 C1178 ( .A(N9), .B(N376), .Z(net500) );
endmodule


module SSTL18DDR3DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   N0, N1, A_, PADN_;
  tri   PAD;
  tri   PADN;
  tri   A;

  GTECH_NOT I_0 ( .A(A), .Z(A_) );
  \**TSGEN**  b1 ( .\function (A), .three_state(N0), .\output (PAD) );
  GTECH_NOT I_1 ( .A(TS), .Z(N0) );
  \**TSGEN**  b2 ( .\function (A_), .three_state(N1), .\output (PADN) );
  GTECH_NOT I_2 ( .A(TS), .Z(N1) );
  GTECH_NOT I_3 ( .A(PADN), .Z(PADN_) );
  GTECH_AND3 a4 ( .A(PAD), .B(PADN_), .C(RI), .Z(Z) );
endmodule


module SSTL18DDR3INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, 
        dq_o, dqs_o, dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_DQ, 
        ts_DQS, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, 
        dq_i, dqs_i, dqsbar_i, dm_i, odt_i, resetbar_i );
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] ba_i;
  input [13:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_DQ, ts_DQS, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i,
         odt_i, resetbar_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad, resetbar_pad;
  wire   ck_o, cke_o, casbar_o, rasbar_o, csbar_o, webar_o, odt_o, resetbar_o;
  wire   [2:0] ba_o;
  wire   [13:0] a_o;
  wire   [1:0] dm_o;
  tri   ck_pad;
  tri   ckbar_pad;
  tri   cke_pad;
  tri   csbar_pad;
  tri   rasbar_pad;
  tri   casbar_pad;
  tri   webar_pad;
  tri   [2:0] ba_pad;
  tri   [13:0] a_pad;
  tri   [1:0] dm_pad;
  tri   odt_pad;
  tri   resetbar_pad;
  tri   [15:0] dq_pad;
  tri   [1:0] dqs_pad;
  tri   [1:0] dqsbar_pad;
  tri   ck_i;
  tri   [15:0] dq_i;
  tri   [1:0] dqs_i;
  tri   [1:0] dm_i;

  SSTL18DDR3DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(ck_o), .A(ck_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_45 cke_sstl ( .PAD(cke_pad), .Z(cke_o), .A(cke_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_44 casbar_sstl ( .PAD(casbar_pad), .Z(casbar_o), .A(casbar_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_43 rasbar_sstl ( .PAD(rasbar_pad), .Z(rasbar_o), .A(rasbar_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_42 csbar_sstl ( .PAD(csbar_pad), .Z(csbar_o), .A(csbar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_41 webar_sstl ( .PAD(webar_pad), .Z(webar_o), .A(webar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_40 odt_sstl ( .PAD(odt_pad), .Z(odt_o), .A(odt_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_39 resetbar_sstl ( .PAD(resetbar_pad), .Z(resetbar_o), .A(
        resetbar_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_38 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(ba_o[0]), .A(ba_i[0]), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_37 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(ba_o[1]), .A(ba_i[1]), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_36 BA_2__sstl_ba ( .PAD(ba_pad[2]), .Z(ba_o[2]), .A(ba_i[2]), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_35 A_0__sstl_a ( .PAD(a_pad[0]), .Z(a_o[0]), .A(a_i[0]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_34 A_1__sstl_a ( .PAD(a_pad[1]), .Z(a_o[1]), .A(a_i[1]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_33 A_2__sstl_a ( .PAD(a_pad[2]), .Z(a_o[2]), .A(a_i[2]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_32 A_3__sstl_a ( .PAD(a_pad[3]), .Z(a_o[3]), .A(a_i[3]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_31 A_4__sstl_a ( .PAD(a_pad[4]), .Z(a_o[4]), .A(a_i[4]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_30 A_5__sstl_a ( .PAD(a_pad[5]), .Z(a_o[5]), .A(a_i[5]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_29 A_6__sstl_a ( .PAD(a_pad[6]), .Z(a_o[6]), .A(a_i[6]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_28 A_7__sstl_a ( .PAD(a_pad[7]), .Z(a_o[7]), .A(a_i[7]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_27 A_8__sstl_a ( .PAD(a_pad[8]), .Z(a_o[8]), .A(a_i[8]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_26 A_9__sstl_a ( .PAD(a_pad[9]), .Z(a_o[9]), .A(a_i[9]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_25 A_10__sstl_a ( .PAD(a_pad[10]), .Z(a_o[10]), .A(a_i[10]), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_24 A_11__sstl_a ( .PAD(a_pad[11]), .Z(a_o[11]), .A(a_i[11]), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_23 A_12__sstl_a ( .PAD(a_pad[12]), .Z(a_o[12]), .A(a_i[12]), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_22 A_13__sstl_a ( .PAD(a_pad[13]), .Z(a_o[13]), .A(a_i[13]), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_DQ) );
  SSTL18DDR3_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_DQS) );
  SSTL18DDR3_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_DQS) );
  SSTL18DDR3_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_DQS) );
  SSTL18DDR3_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_DQS) );
  SSTL18DDR3_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(dm_o[0]), .A(dm_i[0]), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(dm_o[1]), .A(dm_i[1]), .RI(
        1'b0), .TS(1'b1) );
endmodule


module ddr3_controller ( dout, raddr, fillcount, notfull, ready, ck_pad, 
        ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, webar_pad, 
        ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, validout, dq_pad, 
        dqs_pad, dqsbar_pad, clk, reset, read, cmd, din, addr, initddr, sz, op
 );
  output [15:0] dout;
  output [25:0] raddr;
  output [5:0] fillcount;
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [15:0] din;
  input [25:0] addr;
  input [1:0] sz;
  input [2:0] op;
  input clk, reset, read, initddr;
  output notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad,
         casbar_pad, webar_pad, odt_pad, resetbar_pad, validout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, put, N31, N32, N33, N34, IN_empty, IN_full, CMD_full,
         RETURN_empty, init_csbar, init_rasbar, init_casbar, init_webar,
         init_odt, init_ts_con, init_cke, init_resetbar, N35, N36, ts_DQ, N37,
         N38, ts_DQS, N39, N40, N41, N42, N43, N44, csbar_i, N45, N46,
         rasbar_i, N47, N48, casbar_i, N49, N50, webar_i, N51, N52, resetbar_i,
         N53, N54, N55, N56, N57, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;
  wire   [5:0] CMD_fillcount;
  wire   [5:0] RETURN_fillcount;
  wire   [2:0] init_ba;
  wire   [13:0] init_a;
  wire   [13:0] a_i;
  wire   [2:0] ba_i;
  wire   [1:0] dqsbar_i;
  wire   [15:0] dq_o;
  wire   [1:0] dqs_o;
  wire   [1:0] dqsbar_o;
  tri   ready;
  tri   ck_pad;
  tri   ckbar_pad;
  tri   cke_pad;
  tri   csbar_pad;
  tri   rasbar_pad;
  tri   casbar_pad;
  tri   webar_pad;
  tri   [2:0] ba_pad;
  tri   [13:0] a_pad;
  tri   [1:0] dm_pad;
  tri   odt_pad;
  tri   resetbar_pad;
  tri   [15:0] dq_pad;
  tri   [1:0] dqs_pad;
  tri   [1:0] dqsbar_pad;
  tri   clk;
  tri   reset;
  tri   ck_i;
  tri   IN_get;
  tri   [15:0] IN_data_out;
  tri   CMD_get;
  tri   [33:0] CMD_data_out;
  tri   CMD_empty;
  tri   RETURN_put;
  tri   RETURN_full;
  tri   [25:0] RETURN_address;
  tri   [15:0] RETURN_data;
  tri   csbar;
  tri   rasbar;
  tri   casbar;
  tri   webar;
  tri   [2:0] ba;
  tri   [13:0] a;
  tri   [1:0] dm_i;
  tri   [1:0] dqs_i;
  tri   [15:0] dq_i;
  tri   ts_i;
  tri   resetbar;

  GTECH_AND2 C10 ( .A(N23), .B(N24), .Z(N25) );
  GTECH_OR2 C12 ( .A(cmd[1]), .B(N26), .Z(N27) );
  GTECH_OR2 C14 ( .A(N28), .B(cmd[0]), .Z(N29) );
  \**SEQGEN**  ck_i_reg ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ck_i), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  FIFO_DEPTH_P25_WIDTH16 FIFO_IN ( .clk(clk), .reset(reset), .data_in(din), 
        .put(put), .get(IN_get), .data_out(IN_data_out), .empty(IN_empty), 
        .full(IN_full), .fillcount(fillcount) );
  FIFO_DEPTH_P25_WIDTH34 FIFO_CMD ( .clk(clk), .reset(reset), .data_in({cmd, 
        addr, op, sz}), .put(put), .get(CMD_get), .data_out(CMD_data_out), 
        .empty(CMD_empty), .full(CMD_full), .fillcount(CMD_fillcount) );
  FIFO_DEPTH_P25_WIDTH42 FIFO_RETURN ( .clk(clk), .reset(reset), .data_in({
        RETURN_address, RETURN_data}), .put(RETURN_put), .get(read), 
        .data_out({raddr, dout}), .empty(RETURN_empty), .full(RETURN_full), 
        .fillcount(RETURN_fillcount) );
  ddr3_init_engine XINIT ( .ready(ready), .csbar(init_csbar), .rasbar(
        init_rasbar), .casbar(init_casbar), .webar(init_webar), .ba(init_ba), 
        .a(init_a), .dm({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}), 
        .odt(init_odt), .ts_con(init_ts_con), .cke(init_cke), .resetbar(
        init_resetbar), .clk(clk), .reset(reset), .init(initddr), .ck(ck_i) );
  Processing_logic process_logic_ddr3 ( .DATA_get(IN_get), .CMD_get(CMD_get), 
        .RETURN_put(RETURN_put), .RETURN_address(RETURN_address), 
        .RETURN_data(RETURN_data), .cs_bar(csbar), .ras_bar(rasbar), .cas_bar(
        casbar), .we_bar(webar), .BA(ba), .A(a), .DM(dm_i), .DQS_out(dqs_i), 
        .DQ_out(dq_i), .ts_con(ts_i), .resetbar(resetbar), .clk(clk), .ck(ck_i), .reset(reset), .ready(ready), .CMD_empty(CMD_empty), .CMD_data_out(
        CMD_data_out), .DATA_data_out(IN_data_out), .RETURN_full(RETURN_full), 
        .DQS_in(dqs_pad), .DQ_in(dq_pad) );
  SSTL18DDR3INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .resetbar_pad(
        resetbar_pad), .dq_o(dq_o), .dqs_o(dqs_o), .dqsbar_o(dqsbar_o), 
        .dq_pad(dq_pad), .dqs_pad(dqs_pad), .dqsbar_pad(dqsbar_pad), .ri_i(
        1'b1), .ts_DQ(ts_DQ), .ts_DQS(ts_DQS), .ck_i(ck_i), .cke_i(init_cke), 
        .csbar_i(csbar_i), .rasbar_i(rasbar_i), .casbar_i(casbar_i), .webar_i(
        webar_i), .ba_i(ba_i), .a_i(a_i), .dq_i(dq_i), .dqs_i(dqs_i), 
        .dqsbar_i(dqsbar_i), .dm_i(dm_i), .odt_i(init_odt), .resetbar_i(
        resetbar_i) );
  SELECT_OP C106 ( .DATA1(N30), .DATA2(1'b0), .CONTROL1(N0), .CONTROL2(N22), 
        .Z(put) );
  GTECH_BUF B_0 ( .A(N21), .Z(N0) );
  SELECT_OP C107 ( .DATA1(1'b1), .DATA2(N33), .CONTROL1(N1), .CONTROL2(N2), 
        .Z(N34) );
  GTECH_BUF B_1 ( .A(N32), .Z(N1) );
  GTECH_BUF B_2 ( .A(N31), .Z(N2) );
  SELECT_OP C108 ( .DATA1(ts_i), .DATA2(init_ts_con), .CONTROL1(N3), 
        .CONTROL2(N4), .Z(ts_DQ) );
  GTECH_BUF B_3 ( .A(N36), .Z(N3) );
  GTECH_BUF B_4 ( .A(N35), .Z(N4) );
  SELECT_OP C109 ( .DATA1(ts_i), .DATA2(init_ts_con), .CONTROL1(N5), 
        .CONTROL2(N6), .Z(ts_DQS) );
  GTECH_BUF B_5 ( .A(N38), .Z(N5) );
  GTECH_BUF B_6 ( .A(N37), .Z(N6) );
  SELECT_OP C110 ( .DATA1(a), .DATA2(init_a), .CONTROL1(N7), .CONTROL2(N8), 
        .Z(a_i) );
  GTECH_BUF B_7 ( .A(N40), .Z(N7) );
  GTECH_BUF B_8 ( .A(N39), .Z(N8) );
  SELECT_OP C111 ( .DATA1(ba), .DATA2(init_ba), .CONTROL1(N9), .CONTROL2(N10), 
        .Z(ba_i) );
  GTECH_BUF B_9 ( .A(N42), .Z(N9) );
  GTECH_BUF B_10 ( .A(N41), .Z(N10) );
  SELECT_OP C112 ( .DATA1(csbar), .DATA2(init_csbar), .CONTROL1(N11), 
        .CONTROL2(N12), .Z(csbar_i) );
  GTECH_BUF B_11 ( .A(N44), .Z(N11) );
  GTECH_BUF B_12 ( .A(N43), .Z(N12) );
  SELECT_OP C113 ( .DATA1(rasbar), .DATA2(init_rasbar), .CONTROL1(N13), 
        .CONTROL2(N14), .Z(rasbar_i) );
  GTECH_BUF B_13 ( .A(N46), .Z(N13) );
  GTECH_BUF B_14 ( .A(N45), .Z(N14) );
  SELECT_OP C114 ( .DATA1(casbar), .DATA2(init_casbar), .CONTROL1(N15), 
        .CONTROL2(N16), .Z(casbar_i) );
  GTECH_BUF B_15 ( .A(N48), .Z(N15) );
  GTECH_BUF B_16 ( .A(N47), .Z(N16) );
  SELECT_OP C115 ( .DATA1(webar), .DATA2(init_webar), .CONTROL1(N17), 
        .CONTROL2(N18), .Z(webar_i) );
  GTECH_BUF B_17 ( .A(N50), .Z(N17) );
  GTECH_BUF B_18 ( .A(N49), .Z(N18) );
  SELECT_OP C116 ( .DATA1(resetbar), .DATA2(init_resetbar), .CONTROL1(N19), 
        .CONTROL2(N20), .Z(resetbar_i) );
  GTECH_BUF B_19 ( .A(N52), .Z(N19) );
  GTECH_BUF B_20 ( .A(N51), .Z(N20) );
  GTECH_NOT I_0 ( .A(cmd[2]), .Z(N21) );
  GTECH_NOT I_1 ( .A(N21), .Z(N22) );
  GTECH_NOT I_2 ( .A(cmd[1]), .Z(N23) );
  GTECH_NOT I_3 ( .A(cmd[0]), .Z(N24) );
  GTECH_NOT I_4 ( .A(cmd[0]), .Z(N26) );
  GTECH_NOT I_5 ( .A(cmd[1]), .Z(N28) );
  GTECH_OR2 C126 ( .A(N54), .B(N55), .Z(N30) );
  GTECH_OR2 C127 ( .A(N25), .B(N53), .Z(N54) );
  GTECH_NOT I_6 ( .A(N27), .Z(N53) );
  GTECH_NOT I_7 ( .A(N29), .Z(N55) );
  GTECH_NOT I_8 ( .A(reset), .Z(N31) );
  GTECH_BUF B_21 ( .A(reset), .Z(N32) );
  GTECH_NOT I_9 ( .A(ck_i), .Z(N33) );
  GTECH_AND2 C135 ( .A(N56), .B(N57), .Z(notfull) );
  GTECH_NOT I_10 ( .A(CMD_full), .Z(N56) );
  GTECH_NOT I_11 ( .A(IN_full), .Z(N57) );
  GTECH_NOT I_12 ( .A(ready), .Z(N35) );
  GTECH_BUF B_22 ( .A(ready), .Z(N36) );
  GTECH_NOT I_13 ( .A(ready), .Z(N37) );
  GTECH_BUF B_23 ( .A(ready), .Z(N38) );
  GTECH_NOT I_14 ( .A(ready), .Z(N39) );
  GTECH_BUF B_24 ( .A(ready), .Z(N40) );
  GTECH_NOT I_15 ( .A(ready), .Z(N41) );
  GTECH_BUF B_25 ( .A(ready), .Z(N42) );
  GTECH_NOT I_16 ( .A(ready), .Z(N43) );
  GTECH_BUF B_26 ( .A(ready), .Z(N44) );
  GTECH_NOT I_17 ( .A(ready), .Z(N45) );
  GTECH_BUF B_27 ( .A(ready), .Z(N46) );
  GTECH_NOT I_18 ( .A(ready), .Z(N47) );
  GTECH_BUF B_28 ( .A(ready), .Z(N48) );
  GTECH_NOT I_19 ( .A(ready), .Z(N49) );
  GTECH_BUF B_29 ( .A(ready), .Z(N50) );
  GTECH_NOT I_20 ( .A(ready), .Z(N51) );
  GTECH_BUF B_30 ( .A(ready), .Z(N52) );
  GTECH_NOT I_21 ( .A(dqs_i[1]), .Z(dqsbar_i[1]) );
  GTECH_NOT I_22 ( .A(dqs_i[0]), .Z(dqsbar_i[0]) );
  GTECH_NOT I_23 ( .A(RETURN_empty), .Z(validout) );
endmodule


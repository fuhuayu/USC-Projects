
module maze_router_DW01_add_9 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n52, n54, n55, n56, n57, n59, n60, n61, n62, n65,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n81, n82, n83, n84, n85,
         n92, n93, n94, n95, n96, n99, n100, n105, n106, n107, n108, n109,
         n116, n117, n118, n119, n120, n121, n122, n129, n130, n131, n132,
         n138, n139, n140, n143, n144, n145, n146, n151, n152, n153, n154,
         n155, n162, n163, n164, n165, n166, n167, n175, n176, n177, n178,
         n179, n184, n185, n186, n188, n191, n192, n197, n198, n199, n200,
         n201, n206, n207, n208, n209, n210, n219, n223, n225, n226, n227,
         n228, n229, n230, n235, n236, n237, n238, n239, n246, n247, n248,
         n249, n250, n251, n259, n260, n261, n262, n263, n265, n268, n269,
         n270, n272, n275, n276, n280, n281, n282, n283, n284, n285, n290,
         n291, n292, n293, n294, n300, n302, n303, n307, n308, n309, n310,
         n311, n312, n313, n315, n317, n318, n319, n320, n324, n326, n327,
         n328, n329, n330, n331, n335, n337, n338, n339, n340, n345, n346,
         n347, n348, n350, n352, n353, n354, n355, n357, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746;

  XOR2X1 U7 ( .A(n547), .B(n8), .Y(SUM[31]) );
  XOR2X1 U12 ( .A(n546), .B(n619), .Y(SUM[30]) );
  AOI21X1 U13 ( .A(n746), .B(n509), .C(n44), .Y(n42) );
  OAI21X1 U15 ( .A(n649), .B(n719), .C(n590), .Y(n44) );
  AOI21X1 U17 ( .A(n6), .B(n517), .C(n48), .Y(n46) );
  OAI21X1 U19 ( .A(n648), .B(n679), .C(n589), .Y(n48) );
  AOI21X1 U21 ( .A(n728), .B(n65), .C(n52), .Y(n50) );
  XOR2X1 U28 ( .A(n545), .B(n618), .Y(SUM[29]) );
  AOI21X1 U29 ( .A(n746), .B(n508), .C(n57), .Y(n55) );
  OAI21X1 U31 ( .A(n591), .B(n719), .C(n587), .Y(n57) );
  AOI21X1 U33 ( .A(n6), .B(n516), .C(n61), .Y(n59) );
  OAI21X1 U35 ( .A(n672), .B(n678), .C(n655), .Y(n61) );
  XOR2X1 U44 ( .A(n544), .B(n617), .Y(SUM[28]) );
  AOI21X1 U45 ( .A(n746), .B(n507), .C(n70), .Y(n68) );
  OAI21X1 U47 ( .A(n646), .B(n719), .C(n586), .Y(n70) );
  AOI21X1 U49 ( .A(n6), .B(n73), .C(n74), .Y(n72) );
  AOI21X1 U53 ( .A(n740), .B(n566), .C(n567), .Y(n76) );
  XOR2X1 U60 ( .A(n543), .B(n616), .Y(SUM[27]) );
  AOI21X1 U61 ( .A(n746), .B(n506), .C(n83), .Y(n81) );
  OAI21X1 U63 ( .A(n645), .B(n719), .C(n585), .Y(n83) );
  AOI21X1 U65 ( .A(n6), .B(n724), .C(n566), .Y(n85) );
  XOR2X1 U74 ( .A(n542), .B(n615), .Y(SUM[26]) );
  AOI21X1 U75 ( .A(n746), .B(n505), .C(n94), .Y(n92) );
  OAI21X1 U77 ( .A(n95), .B(n719), .C(n96), .Y(n94) );
  OAI21X1 U81 ( .A(n592), .B(n667), .C(n584), .Y(n6) );
  AOI21X1 U83 ( .A(n737), .B(n564), .C(n565), .Y(n100) );
  XOR2X1 U90 ( .A(n541), .B(n614), .Y(SUM[25]) );
  AOI21X1 U91 ( .A(n746), .B(n504), .C(n107), .Y(n105) );
  OAI21X1 U93 ( .A(n515), .B(n719), .C(n582), .Y(n107) );
  AOI21X1 U95 ( .A(n122), .B(n726), .C(n564), .Y(n109) );
  XOR2X1 U104 ( .A(n540), .B(n613), .Y(SUM[24]) );
  AOI21X1 U105 ( .A(n746), .B(n503), .C(n118), .Y(n116) );
  OAI21X1 U107 ( .A(n685), .B(n719), .C(n668), .Y(n118) );
  AOI21X1 U113 ( .A(n734), .B(n562), .C(n563), .Y(n120) );
  XOR2X1 U120 ( .A(n539), .B(n612), .Y(SUM[23]) );
  AOI21X1 U121 ( .A(n746), .B(n595), .C(n131), .Y(n129) );
  OAI21X1 U123 ( .A(n671), .B(n719), .C(n654), .Y(n131) );
  XOR2X1 U132 ( .A(n597), .B(n611), .Y(SUM[22]) );
  AOI21X1 U133 ( .A(n746), .B(n139), .C(n140), .Y(n138) );
  AOI21X1 U137 ( .A(n186), .B(n594), .C(n144), .Y(n4) );
  OAI21X1 U139 ( .A(n644), .B(n665), .C(n720), .Y(n144) );
  AOI21X1 U141 ( .A(n741), .B(n560), .C(n561), .Y(n146) );
  XOR2X1 U148 ( .A(n538), .B(n610), .Y(SUM[21]) );
  AOI21X1 U149 ( .A(n745), .B(n502), .C(n153), .Y(n151) );
  OAI21X1 U151 ( .A(n642), .B(n188), .C(n581), .Y(n153) );
  AOI21X1 U153 ( .A(n664), .B(n725), .C(n560), .Y(n155) );
  XOR2X1 U162 ( .A(n537), .B(n609), .Y(SUM[20]) );
  AOI21X1 U163 ( .A(n745), .B(n501), .C(n164), .Y(n162) );
  OAI21X1 U165 ( .A(n683), .B(n188), .C(n665), .Y(n164) );
  AOI21X1 U171 ( .A(n733), .B(n179), .C(n559), .Y(n166) );
  XOR2X1 U178 ( .A(n536), .B(n699), .Y(SUM[19]) );
  AOI21X1 U179 ( .A(n745), .B(n500), .C(n177), .Y(n175) );
  OAI21X1 U181 ( .A(n710), .B(n188), .C(n707), .Y(n177) );
  XOR2X1 U190 ( .A(n535), .B(n608), .Y(SUM[18]) );
  AOI21X1 U191 ( .A(n745), .B(n659), .C(n186), .Y(n184) );
  OAI21X1 U197 ( .A(n641), .B(n675), .C(n579), .Y(n186) );
  AOI21X1 U199 ( .A(n735), .B(n201), .C(n558), .Y(n192) );
  XOR2X1 U206 ( .A(n534), .B(n607), .Y(SUM[17]) );
  AOI21X1 U207 ( .A(n745), .B(n499), .C(n199), .Y(n197) );
  OAI21X1 U209 ( .A(n670), .B(n676), .C(n653), .Y(n199) );
  XOR2X1 U218 ( .A(n533), .B(n606), .Y(SUM[16]) );
  AOI21X1 U219 ( .A(n745), .B(n207), .C(n208), .Y(n206) );
  AOI21X1 U227 ( .A(n743), .B(n223), .C(n557), .Y(n210) );
  XNOR2X1 U234 ( .A(n745), .B(n716), .Y(SUM[15]) );
  AOI21X1 U235 ( .A(n745), .B(n730), .C(n223), .Y(n219) );
  XOR2X1 U242 ( .A(n532), .B(n605), .Y(SUM[14]) );
  OAI21X1 U243 ( .A(n514), .B(n522), .C(n519), .Y(n3) );
  AOI21X1 U245 ( .A(n270), .B(n513), .C(n228), .Y(n226) );
  OAI21X1 U247 ( .A(n640), .B(n663), .C(n577), .Y(n228) );
  AOI21X1 U249 ( .A(n742), .B(n555), .C(n556), .Y(n230) );
  XOR2X1 U256 ( .A(n531), .B(n604), .Y(SUM[13]) );
  AOI21X1 U257 ( .A(n308), .B(n498), .C(n237), .Y(n235) );
  OAI21X1 U259 ( .A(n639), .B(n272), .C(n575), .Y(n237) );
  AOI21X1 U261 ( .A(n662), .B(n727), .C(n555), .Y(n239) );
  XOR2X1 U270 ( .A(n530), .B(n603), .Y(SUM[12]) );
  AOI21X1 U271 ( .A(n308), .B(n497), .C(n248), .Y(n246) );
  OAI21X1 U273 ( .A(n681), .B(n272), .C(n663), .Y(n248) );
  AOI21X1 U279 ( .A(n732), .B(n265), .C(n554), .Y(n250) );
  XOR2X1 U286 ( .A(n529), .B(n602), .Y(SUM[11]) );
  AOI21X1 U287 ( .A(n308), .B(n496), .C(n261), .Y(n259) );
  OAI21X1 U289 ( .A(n709), .B(n272), .C(n701), .Y(n261) );
  XOR2X1 U298 ( .A(n528), .B(n601), .Y(SUM[10]) );
  AOI21X1 U299 ( .A(n308), .B(n661), .C(n270), .Y(n268) );
  OAI21X1 U305 ( .A(n638), .B(n523), .C(n574), .Y(n270) );
  AOI21X1 U307 ( .A(n731), .B(n285), .C(n280), .Y(n276) );
  XOR2X1 U314 ( .A(n527), .B(n600), .Y(SUM[9]) );
  AOI21X1 U315 ( .A(n308), .B(n495), .C(n283), .Y(n281) );
  OAI21X1 U317 ( .A(n669), .B(n673), .C(n652), .Y(n283) );
  XOR2X1 U326 ( .A(n526), .B(n599), .Y(SUM[8]) );
  AOI21X1 U327 ( .A(n308), .B(n291), .C(n292), .Y(n290) );
  AOI21X1 U335 ( .A(n738), .B(n307), .C(n300), .Y(n294) );
  XNOR2X1 U342 ( .A(n308), .B(n714), .Y(SUM[7]) );
  AOI21X1 U343 ( .A(n308), .B(n736), .C(n307), .Y(n303) );
  XNOR2X1 U350 ( .A(n318), .B(n713), .Y(SUM[6]) );
  AOI21X1 U352 ( .A(n346), .B(n510), .C(n311), .Y(n309) );
  OAI21X1 U354 ( .A(n637), .B(n708), .C(n572), .Y(n311) );
  AOI21X1 U356 ( .A(n744), .B(n324), .C(n315), .Y(n313) );
  XNOR2X1 U363 ( .A(n327), .B(n717), .Y(SUM[5]) );
  OAI21X1 U364 ( .A(n520), .B(n345), .C(n518), .Y(n318) );
  AOI21X1 U366 ( .A(n331), .B(n723), .C(n324), .Y(n320) );
  XNOR2X1 U375 ( .A(n338), .B(n712), .Y(SUM[4]) );
  OAI21X1 U376 ( .A(n551), .B(n345), .C(n708), .Y(n327) );
  AOI21X1 U382 ( .A(n739), .B(n340), .C(n335), .Y(n329) );
  XOR2X1 U389 ( .A(n345), .B(n696), .Y(SUM[3]) );
  OAI21X1 U390 ( .A(n700), .B(n345), .C(n718), .Y(n338) );
  XNOR2X1 U399 ( .A(n353), .B(n715), .Y(SUM[2]) );
  OAI21X1 U401 ( .A(n596), .B(n688), .C(n571), .Y(n346) );
  AOI21X1 U403 ( .A(n729), .B(n357), .C(n350), .Y(n348) );
  XOR2X1 U410 ( .A(n690), .B(n598), .Y(SUM[1]) );
  OAI21X1 U411 ( .A(n636), .B(n689), .C(n651), .Y(n353) );
  OR2X2 U428 ( .A(A[24]), .B(B[24]), .Y(n734) );
  AND2X1 U429 ( .A(n729), .B(n354), .Y(n347) );
  BUFX2 U430 ( .A(n3), .Y(n745) );
  OR2X2 U431 ( .A(A[20]), .B(B[20]), .Y(n733) );
  OR2X2 U432 ( .A(n550), .B(n669), .Y(n282) );
  INVX1 U433 ( .A(n282), .Y(n495) );
  OR2X2 U434 ( .A(n660), .B(n709), .Y(n260) );
  INVX1 U435 ( .A(n260), .Y(n496) );
  OR2X2 U436 ( .A(n660), .B(n681), .Y(n247) );
  INVX1 U437 ( .A(n247), .Y(n497) );
  OR2X2 U438 ( .A(n660), .B(n639), .Y(n236) );
  INVX1 U439 ( .A(n236), .Y(n498) );
  OR2X2 U440 ( .A(n657), .B(n670), .Y(n198) );
  INVX1 U441 ( .A(n198), .Y(n499) );
  OR2X2 U442 ( .A(n185), .B(n710), .Y(n176) );
  INVX1 U443 ( .A(n176), .Y(n500) );
  OR2X2 U444 ( .A(n185), .B(n683), .Y(n163) );
  INVX1 U445 ( .A(n163), .Y(n501) );
  OR2X2 U446 ( .A(n185), .B(n643), .Y(n152) );
  INVX1 U447 ( .A(n152), .Y(n502) );
  OR2X2 U448 ( .A(n692), .B(n685), .Y(n117) );
  INVX1 U449 ( .A(n117), .Y(n503) );
  OR2X2 U450 ( .A(n691), .B(n515), .Y(n106) );
  INVX1 U451 ( .A(n106), .Y(n504) );
  OR2X2 U452 ( .A(n691), .B(n95), .Y(n93) );
  INVX1 U453 ( .A(n93), .Y(n505) );
  OR2X2 U454 ( .A(n693), .B(n645), .Y(n82) );
  INVX1 U455 ( .A(n82), .Y(n506) );
  OR2X2 U456 ( .A(n692), .B(n646), .Y(n69) );
  INVX1 U457 ( .A(n69), .Y(n507) );
  OR2X2 U458 ( .A(n693), .B(n591), .Y(n56) );
  INVX1 U459 ( .A(n56), .Y(n508) );
  OR2X2 U460 ( .A(n692), .B(n649), .Y(n43) );
  INVX1 U461 ( .A(n43), .Y(n509) );
  AND2X2 U462 ( .A(n689), .B(n722), .Y(SUM[0]) );
  AND2X2 U463 ( .A(A[1]), .B(B[1]), .Y(n355) );
  OR2X2 U464 ( .A(B[1]), .B(A[1]), .Y(n354) );
  OR2X2 U465 ( .A(n552), .B(n637), .Y(n310) );
  INVX1 U466 ( .A(n310), .Y(n510) );
  AND2X2 U467 ( .A(B[9]), .B(A[9]), .Y(n285) );
  OR2X2 U468 ( .A(A[9]), .B(B[9]), .Y(n284) );
  AND2X2 U469 ( .A(B[10]), .B(A[10]), .Y(n280) );
  INVX1 U470 ( .A(n280), .Y(n511) );
  AND2X2 U471 ( .A(n731), .B(n284), .Y(n275) );
  OR2X2 U472 ( .A(n549), .B(n570), .Y(n269) );
  INVX1 U473 ( .A(n269), .Y(n512) );
  OR2X2 U474 ( .A(n682), .B(n640), .Y(n227) );
  INVX1 U475 ( .A(n227), .Y(n513) );
  AND2X2 U476 ( .A(n513), .B(n512), .Y(n225) );
  INVX1 U477 ( .A(n225), .Y(n514) );
  OR2X2 U478 ( .A(A[17]), .B(B[17]), .Y(n200) );
  OR2X2 U479 ( .A(n683), .B(n644), .Y(n143) );
  AND2X2 U480 ( .A(n726), .B(n121), .Y(n108) );
  INVX1 U481 ( .A(n108), .Y(n515) );
  OR2X2 U482 ( .A(n658), .B(n672), .Y(n60) );
  INVX1 U483 ( .A(n60), .Y(n516) );
  OR2X2 U484 ( .A(n658), .B(n647), .Y(n47) );
  INVX1 U485 ( .A(n47), .Y(n517) );
  BUFX2 U486 ( .A(n320), .Y(n518) );
  BUFX2 U487 ( .A(n226), .Y(n519) );
  AND2X2 U488 ( .A(n723), .B(n330), .Y(n319) );
  INVX1 U489 ( .A(n319), .Y(n520) );
  OR2X2 U490 ( .A(n656), .B(n641), .Y(n185) );
  INVX1 U491 ( .A(n185), .Y(n521) );
  BUFX2 U492 ( .A(n309), .Y(n522) );
  BUFX2 U493 ( .A(n294), .Y(n523) );
  OR2X2 U494 ( .A(n684), .B(n592), .Y(n7) );
  INVX1 U495 ( .A(n7), .Y(n524) );
  INVX1 U496 ( .A(n7), .Y(n525) );
  BUFX2 U497 ( .A(n303), .Y(n526) );
  BUFX2 U498 ( .A(n290), .Y(n527) );
  BUFX2 U499 ( .A(n281), .Y(n528) );
  BUFX2 U500 ( .A(n268), .Y(n529) );
  BUFX2 U501 ( .A(n259), .Y(n530) );
  BUFX2 U502 ( .A(n246), .Y(n531) );
  BUFX2 U503 ( .A(n235), .Y(n532) );
  BUFX2 U504 ( .A(n219), .Y(n533) );
  BUFX2 U505 ( .A(n206), .Y(n534) );
  BUFX2 U506 ( .A(n197), .Y(n535) );
  BUFX2 U507 ( .A(n184), .Y(n536) );
  BUFX2 U508 ( .A(n175), .Y(n537) );
  BUFX2 U509 ( .A(n162), .Y(n538) );
  BUFX2 U510 ( .A(n138), .Y(n539) );
  BUFX2 U511 ( .A(n129), .Y(n540) );
  BUFX2 U512 ( .A(n116), .Y(n541) );
  BUFX2 U513 ( .A(n105), .Y(n542) );
  BUFX2 U514 ( .A(n92), .Y(n543) );
  BUFX2 U515 ( .A(n81), .Y(n544) );
  BUFX2 U516 ( .A(n68), .Y(n545) );
  BUFX2 U517 ( .A(n55), .Y(n546) );
  BUFX2 U518 ( .A(n42), .Y(n547) );
  AND2X2 U519 ( .A(n738), .B(n736), .Y(n293) );
  INVX1 U520 ( .A(n293), .Y(n548) );
  INVX1 U521 ( .A(n293), .Y(n549) );
  INVX1 U522 ( .A(n293), .Y(n550) );
  AND2X2 U523 ( .A(n739), .B(n339), .Y(n328) );
  INVX1 U524 ( .A(n328), .Y(n551) );
  INVX1 U525 ( .A(n328), .Y(n552) );
  INVX1 U526 ( .A(n328), .Y(n553) );
  AND2X2 U527 ( .A(B[12]), .B(A[12]), .Y(n554) );
  AND2X2 U528 ( .A(B[13]), .B(A[13]), .Y(n555) );
  AND2X2 U529 ( .A(B[14]), .B(A[14]), .Y(n556) );
  AND2X2 U530 ( .A(B[16]), .B(A[16]), .Y(n557) );
  AND2X2 U531 ( .A(B[18]), .B(A[18]), .Y(n558) );
  AND2X2 U532 ( .A(B[20]), .B(A[20]), .Y(n559) );
  AND2X2 U533 ( .A(B[21]), .B(A[21]), .Y(n560) );
  AND2X2 U534 ( .A(B[22]), .B(A[22]), .Y(n561) );
  AND2X2 U535 ( .A(B[23]), .B(A[23]), .Y(n562) );
  AND2X2 U536 ( .A(B[24]), .B(A[24]), .Y(n563) );
  AND2X2 U537 ( .A(B[25]), .B(A[25]), .Y(n564) );
  AND2X2 U538 ( .A(B[26]), .B(A[26]), .Y(n565) );
  AND2X2 U539 ( .A(B[27]), .B(A[27]), .Y(n566) );
  AND2X2 U540 ( .A(B[28]), .B(A[28]), .Y(n567) );
  AND2X2 U541 ( .A(B[29]), .B(A[29]), .Y(n568) );
  AND2X2 U542 ( .A(n516), .B(n525), .Y(n569) );
  INVX1 U543 ( .A(n275), .Y(n570) );
  BUFX2 U544 ( .A(n348), .Y(n571) );
  BUFX2 U545 ( .A(n313), .Y(n572) );
  INVX1 U546 ( .A(n276), .Y(n573) );
  INVX1 U547 ( .A(n573), .Y(n574) );
  BUFX2 U548 ( .A(n239), .Y(n575) );
  INVX1 U549 ( .A(n230), .Y(n576) );
  INVX1 U550 ( .A(n576), .Y(n577) );
  INVX1 U551 ( .A(n192), .Y(n578) );
  INVX1 U552 ( .A(n578), .Y(n579) );
  INVX1 U553 ( .A(n155), .Y(n580) );
  INVX1 U554 ( .A(n580), .Y(n581) );
  BUFX2 U555 ( .A(n109), .Y(n582) );
  INVX1 U556 ( .A(n100), .Y(n583) );
  INVX1 U557 ( .A(n583), .Y(n584) );
  BUFX2 U558 ( .A(n85), .Y(n585) );
  BUFX2 U559 ( .A(n72), .Y(n586) );
  BUFX2 U560 ( .A(n59), .Y(n587) );
  INVX1 U561 ( .A(n50), .Y(n588) );
  INVX1 U562 ( .A(n588), .Y(n589) );
  BUFX2 U563 ( .A(n46), .Y(n590) );
  INVX1 U564 ( .A(n569), .Y(n591) );
  AND2X2 U565 ( .A(n737), .B(n726), .Y(n99) );
  INVX1 U566 ( .A(n99), .Y(n592) );
  OR2X2 U567 ( .A(A[25]), .B(B[25]), .Y(n726) );
  INVX1 U568 ( .A(n143), .Y(n593) );
  INVX1 U569 ( .A(n143), .Y(n594) );
  OR2X2 U570 ( .A(n691), .B(n671), .Y(n130) );
  INVX1 U571 ( .A(n130), .Y(n595) );
  INVX1 U572 ( .A(n347), .Y(n596) );
  BUFX2 U573 ( .A(n151), .Y(n597) );
  AND2X2 U574 ( .A(n651), .B(n354), .Y(n38) );
  INVX1 U575 ( .A(n38), .Y(n598) );
  AND2X2 U576 ( .A(n621), .B(n738), .Y(n31) );
  INVX1 U577 ( .A(n31), .Y(n599) );
  AND2X2 U578 ( .A(n652), .B(n284), .Y(n30) );
  INVX1 U579 ( .A(n30), .Y(n600) );
  AND2X2 U580 ( .A(n511), .B(n731), .Y(n29) );
  INVX1 U581 ( .A(n29), .Y(n601) );
  AND2X2 U582 ( .A(n701), .B(n262), .Y(n28) );
  INVX1 U583 ( .A(n28), .Y(n602) );
  AND2X2 U584 ( .A(n622), .B(n732), .Y(n27) );
  INVX1 U585 ( .A(n27), .Y(n603) );
  AND2X2 U586 ( .A(n623), .B(n727), .Y(n26) );
  INVX1 U587 ( .A(n26), .Y(n604) );
  AND2X2 U588 ( .A(n624), .B(n742), .Y(n25) );
  INVX1 U589 ( .A(n25), .Y(n605) );
  AND2X2 U590 ( .A(n625), .B(n743), .Y(n23) );
  INVX1 U591 ( .A(n23), .Y(n606) );
  AND2X2 U592 ( .A(n653), .B(n200), .Y(n22) );
  INVX1 U593 ( .A(n22), .Y(n607) );
  AND2X2 U594 ( .A(n626), .B(n735), .Y(n21) );
  INVX1 U595 ( .A(n21), .Y(n608) );
  AND2X2 U596 ( .A(n627), .B(n733), .Y(n19) );
  INVX1 U597 ( .A(n19), .Y(n609) );
  AND2X2 U598 ( .A(n628), .B(n725), .Y(n18) );
  INVX1 U599 ( .A(n18), .Y(n610) );
  AND2X2 U600 ( .A(n629), .B(n741), .Y(n17) );
  INVX1 U601 ( .A(n17), .Y(n611) );
  AND2X2 U602 ( .A(n654), .B(n132), .Y(n16) );
  INVX1 U603 ( .A(n16), .Y(n612) );
  AND2X2 U604 ( .A(n630), .B(n734), .Y(n15) );
  INVX1 U605 ( .A(n15), .Y(n613) );
  AND2X2 U606 ( .A(n631), .B(n726), .Y(n14) );
  INVX1 U607 ( .A(n14), .Y(n614) );
  AND2X2 U608 ( .A(n632), .B(n737), .Y(n13) );
  INVX1 U609 ( .A(n13), .Y(n615) );
  AND2X2 U610 ( .A(n633), .B(n724), .Y(n12) );
  INVX1 U611 ( .A(n12), .Y(n616) );
  AND2X2 U612 ( .A(n634), .B(n740), .Y(n11) );
  INVX1 U613 ( .A(n11), .Y(n617) );
  AND2X2 U614 ( .A(n655), .B(n62), .Y(n10) );
  INVX1 U615 ( .A(n10), .Y(n618) );
  AND2X2 U616 ( .A(n635), .B(n728), .Y(n9) );
  INVX1 U617 ( .A(n9), .Y(n619) );
  AND2X2 U618 ( .A(B[8]), .B(A[8]), .Y(n302) );
  INVX1 U619 ( .A(n302), .Y(n620) );
  INVX1 U620 ( .A(n302), .Y(n621) );
  INVX1 U621 ( .A(n554), .Y(n622) );
  INVX1 U622 ( .A(n555), .Y(n623) );
  INVX1 U623 ( .A(n556), .Y(n624) );
  INVX1 U624 ( .A(n557), .Y(n625) );
  INVX1 U625 ( .A(n558), .Y(n626) );
  INVX1 U626 ( .A(n559), .Y(n627) );
  INVX1 U627 ( .A(n560), .Y(n628) );
  INVX1 U628 ( .A(n561), .Y(n629) );
  INVX1 U629 ( .A(n563), .Y(n630) );
  INVX1 U630 ( .A(n564), .Y(n631) );
  INVX1 U631 ( .A(n565), .Y(n632) );
  INVX1 U632 ( .A(n566), .Y(n633) );
  INVX1 U633 ( .A(n567), .Y(n634) );
  AND2X2 U634 ( .A(A[30]), .B(B[30]), .Y(n54) );
  INVX1 U635 ( .A(n54), .Y(n635) );
  INVX1 U636 ( .A(n354), .Y(n636) );
  AND2X2 U637 ( .A(n744), .B(n723), .Y(n312) );
  INVX1 U638 ( .A(n312), .Y(n637) );
  INVX1 U639 ( .A(n275), .Y(n638) );
  OR2X2 U640 ( .A(A[10]), .B(B[10]), .Y(n731) );
  AND2X2 U641 ( .A(n727), .B(n251), .Y(n238) );
  INVX1 U642 ( .A(n238), .Y(n639) );
  AND2X2 U643 ( .A(n742), .B(n727), .Y(n229) );
  INVX1 U644 ( .A(n229), .Y(n640) );
  OR2X2 U645 ( .A(A[13]), .B(B[13]), .Y(n727) );
  AND2X2 U646 ( .A(n735), .B(n200), .Y(n191) );
  INVX1 U647 ( .A(n191), .Y(n641) );
  OR2X2 U648 ( .A(A[18]), .B(B[18]), .Y(n735) );
  AND2X2 U649 ( .A(n725), .B(n167), .Y(n154) );
  INVX1 U650 ( .A(n154), .Y(n642) );
  INVX1 U651 ( .A(n154), .Y(n643) );
  AND2X2 U652 ( .A(n741), .B(n725), .Y(n145) );
  INVX1 U653 ( .A(n145), .Y(n644) );
  AND2X2 U654 ( .A(n724), .B(n524), .Y(n84) );
  INVX1 U655 ( .A(n84), .Y(n645) );
  AND2X2 U656 ( .A(n73), .B(n687), .Y(n71) );
  INVX1 U657 ( .A(n71), .Y(n646) );
  AND2X2 U658 ( .A(n728), .B(n62), .Y(n49) );
  INVX1 U659 ( .A(n49), .Y(n647) );
  INVX1 U660 ( .A(n49), .Y(n648) );
  AND2X2 U661 ( .A(n517), .B(n687), .Y(n45) );
  INVX1 U662 ( .A(n45), .Y(n649) );
  INVX1 U663 ( .A(n355), .Y(n650) );
  INVX1 U664 ( .A(n355), .Y(n651) );
  INVX1 U665 ( .A(n285), .Y(n652) );
  INVX1 U666 ( .A(n201), .Y(n653) );
  AND2X2 U667 ( .A(B[17]), .B(A[17]), .Y(n201) );
  INVX1 U668 ( .A(n562), .Y(n654) );
  INVX1 U669 ( .A(n568), .Y(n655) );
  INVX1 U670 ( .A(n209), .Y(n656) );
  INVX1 U671 ( .A(n209), .Y(n657) );
  AND2X2 U672 ( .A(n743), .B(n730), .Y(n209) );
  INVX1 U673 ( .A(n75), .Y(n658) );
  AND2X2 U674 ( .A(n740), .B(n724), .Y(n75) );
  INVX1 U675 ( .A(n185), .Y(n659) );
  INVX1 U676 ( .A(n512), .Y(n660) );
  INVX1 U677 ( .A(n660), .Y(n661) );
  INVX1 U678 ( .A(n250), .Y(n662) );
  INVX1 U679 ( .A(n662), .Y(n663) );
  INVX1 U680 ( .A(n166), .Y(n664) );
  INVX1 U681 ( .A(n664), .Y(n665) );
  INVX1 U682 ( .A(n120), .Y(n666) );
  INVX1 U683 ( .A(n666), .Y(n667) );
  INVX1 U684 ( .A(n666), .Y(n668) );
  INVX1 U685 ( .A(n284), .Y(n669) );
  INVX1 U686 ( .A(n200), .Y(n670) );
  INVX1 U687 ( .A(n132), .Y(n671) );
  OR2X2 U688 ( .A(A[23]), .B(B[23]), .Y(n132) );
  INVX1 U689 ( .A(n62), .Y(n672) );
  OR2X2 U690 ( .A(A[29]), .B(B[29]), .Y(n62) );
  INVX1 U691 ( .A(n292), .Y(n673) );
  INVX1 U692 ( .A(n210), .Y(n674) );
  INVX1 U693 ( .A(n674), .Y(n675) );
  INVX1 U694 ( .A(n674), .Y(n676) );
  INVX1 U695 ( .A(n76), .Y(n677) );
  INVX1 U696 ( .A(n677), .Y(n678) );
  INVX1 U697 ( .A(n677), .Y(n679) );
  INVX1 U698 ( .A(n682), .Y(n680) );
  INVX1 U699 ( .A(n680), .Y(n681) );
  AND2X2 U700 ( .A(n732), .B(n262), .Y(n249) );
  INVX1 U701 ( .A(n249), .Y(n682) );
  AND2X2 U702 ( .A(n733), .B(n178), .Y(n165) );
  INVX1 U703 ( .A(n165), .Y(n683) );
  INVX1 U704 ( .A(n119), .Y(n684) );
  INVX1 U705 ( .A(n119), .Y(n685) );
  AND2X2 U706 ( .A(n734), .B(n132), .Y(n119) );
  INVX1 U707 ( .A(n525), .Y(n686) );
  INVX1 U708 ( .A(n686), .Y(n687) );
  INVX1 U709 ( .A(n1), .Y(n688) );
  INVX1 U710 ( .A(n1), .Y(n689) );
  INVX1 U711 ( .A(n1), .Y(n690) );
  AND2X2 U712 ( .A(B[0]), .B(A[0]), .Y(n1) );
  INVX1 U713 ( .A(n5), .Y(n691) );
  INVX1 U714 ( .A(n5), .Y(n692) );
  INVX1 U715 ( .A(n5), .Y(n693) );
  AND2X2 U716 ( .A(n593), .B(n521), .Y(n5) );
  OR2X2 U717 ( .A(A[26]), .B(B[26]), .Y(n737) );
  OR2X2 U718 ( .A(A[27]), .B(B[27]), .Y(n724) );
  OR2X2 U719 ( .A(A[14]), .B(B[14]), .Y(n742) );
  OR2X2 U720 ( .A(A[0]), .B(B[0]), .Y(n722) );
  OR2X2 U721 ( .A(A[16]), .B(B[16]), .Y(n743) );
  OR2X2 U722 ( .A(A[28]), .B(B[28]), .Y(n740) );
  OR2X2 U723 ( .A(A[21]), .B(B[21]), .Y(n725) );
  OR2X2 U724 ( .A(A[8]), .B(B[8]), .Y(n738) );
  AND2X2 U725 ( .A(A[2]), .B(B[2]), .Y(n352) );
  INVX1 U726 ( .A(n352), .Y(n694) );
  INVX1 U727 ( .A(n352), .Y(n695) );
  AND2X2 U728 ( .A(n718), .B(n339), .Y(n36) );
  INVX1 U729 ( .A(n36), .Y(n696) );
  AND2X2 U730 ( .A(B[4]), .B(A[4]), .Y(n337) );
  INVX1 U731 ( .A(n337), .Y(n697) );
  INVX1 U732 ( .A(n337), .Y(n698) );
  AND2X2 U733 ( .A(n707), .B(n178), .Y(n20) );
  INVX1 U734 ( .A(n20), .Y(n699) );
  OR2X2 U735 ( .A(A[3]), .B(B[3]), .Y(n339) );
  INVX1 U736 ( .A(n339), .Y(n700) );
  AND2X2 U737 ( .A(B[11]), .B(A[11]), .Y(n263) );
  INVX1 U738 ( .A(n263), .Y(n701) );
  AND2X2 U739 ( .A(B[15]), .B(A[15]), .Y(n223) );
  INVX1 U740 ( .A(n223), .Y(n702) );
  AND2X2 U741 ( .A(B[7]), .B(A[7]), .Y(n307) );
  INVX1 U742 ( .A(n307), .Y(n703) );
  AND2X2 U743 ( .A(B[6]), .B(A[6]), .Y(n317) );
  INVX1 U744 ( .A(n317), .Y(n704) );
  AND2X2 U745 ( .A(A[5]), .B(B[5]), .Y(n326) );
  INVX1 U746 ( .A(n326), .Y(n705) );
  INVX1 U747 ( .A(n326), .Y(n706) );
  AND2X2 U748 ( .A(B[19]), .B(A[19]), .Y(n179) );
  INVX1 U749 ( .A(n179), .Y(n707) );
  BUFX2 U750 ( .A(n329), .Y(n708) );
  OR2X2 U751 ( .A(A[11]), .B(B[11]), .Y(n262) );
  INVX1 U752 ( .A(n262), .Y(n709) );
  OR2X2 U753 ( .A(A[19]), .B(B[19]), .Y(n178) );
  INVX1 U754 ( .A(n178), .Y(n710) );
  OR2X2 U755 ( .A(B[31]), .B(A[31]), .Y(n40) );
  INVX1 U756 ( .A(n40), .Y(n711) );
  OR2X2 U757 ( .A(n721), .B(n711), .Y(n8) );
  AND2X2 U758 ( .A(n698), .B(n739), .Y(n35) );
  INVX1 U759 ( .A(n35), .Y(n712) );
  OR2X2 U760 ( .A(A[4]), .B(B[4]), .Y(n739) );
  AND2X2 U761 ( .A(n704), .B(n744), .Y(n33) );
  INVX1 U762 ( .A(n33), .Y(n713) );
  OR2X2 U763 ( .A(A[6]), .B(B[6]), .Y(n744) );
  AND2X2 U764 ( .A(n703), .B(n736), .Y(n32) );
  INVX1 U765 ( .A(n32), .Y(n714) );
  OR2X2 U766 ( .A(A[7]), .B(B[7]), .Y(n736) );
  AND2X2 U767 ( .A(n695), .B(n729), .Y(n37) );
  INVX1 U768 ( .A(n37), .Y(n715) );
  OR2X2 U769 ( .A(B[2]), .B(A[2]), .Y(n729) );
  AND2X2 U770 ( .A(n702), .B(n730), .Y(n24) );
  INVX1 U771 ( .A(n24), .Y(n716) );
  OR2X2 U772 ( .A(A[15]), .B(B[15]), .Y(n730) );
  AND2X2 U773 ( .A(n706), .B(n723), .Y(n34) );
  INVX1 U774 ( .A(n34), .Y(n717) );
  OR2X2 U775 ( .A(B[5]), .B(A[5]), .Y(n723) );
  AND2X2 U776 ( .A(B[3]), .B(A[3]), .Y(n340) );
  INVX1 U777 ( .A(n340), .Y(n718) );
  BUFX2 U778 ( .A(n4), .Y(n719) );
  BUFX2 U779 ( .A(n146), .Y(n720) );
  OR2X2 U780 ( .A(A[22]), .B(B[22]), .Y(n741) );
  BUFX2 U781 ( .A(n3), .Y(n746) );
  INVX1 U782 ( .A(n522), .Y(n308) );
  INVX1 U783 ( .A(n548), .Y(n291) );
  INVX1 U784 ( .A(n523), .Y(n292) );
  INVX1 U785 ( .A(n525), .Y(n95) );
  INVX1 U786 ( .A(n693), .Y(n139) );
  INVX1 U787 ( .A(n719), .Y(n140) );
  INVX1 U788 ( .A(n657), .Y(n207) );
  INVX1 U789 ( .A(n676), .Y(n208) );
  INVX1 U790 ( .A(n6), .Y(n96) );
  INVX1 U791 ( .A(n346), .Y(n345) );
  INVX1 U792 ( .A(n186), .Y(n188) );
  INVX1 U793 ( .A(n270), .Y(n272) );
  INVX1 U794 ( .A(n679), .Y(n74) );
  INVX1 U795 ( .A(n681), .Y(n251) );
  INVX1 U796 ( .A(n684), .Y(n121) );
  INVX1 U797 ( .A(n683), .Y(n167) );
  INVX1 U798 ( .A(n658), .Y(n73) );
  INVX1 U799 ( .A(n708), .Y(n331) );
  INVX1 U800 ( .A(n620), .Y(n300) );
  INVX1 U801 ( .A(n694), .Y(n350) );
  INVX1 U802 ( .A(n553), .Y(n330) );
  INVX1 U803 ( .A(n701), .Y(n265) );
  INVX1 U804 ( .A(n697), .Y(n335) );
  INVX1 U805 ( .A(n635), .Y(n52) );
  INVX1 U806 ( .A(n668), .Y(n122) );
  INVX1 U807 ( .A(n655), .Y(n65) );
  INVX1 U808 ( .A(n650), .Y(n357) );
  INVX1 U809 ( .A(n705), .Y(n324) );
  INVX1 U810 ( .A(n704), .Y(n315) );
  AND2X1 U811 ( .A(A[31]), .B(B[31]), .Y(n721) );
  OR2X1 U812 ( .A(B[30]), .B(A[30]), .Y(n728) );
  OR2X1 U813 ( .A(A[12]), .B(B[12]), .Y(n732) );
endmodule


module maze_router_DW_mult_tc_2 ( a, b, product );
  input [31:0] a;
  input [3:0] b;
  output [35:0] product;
  wire   n1, n2, n3, n7, n9, n11, n12, n13, n16, n17, n19, n20, n21, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n36, n37, n38, n39, n40, n41,
         n43, n45, n47, n49, n50, n51, n52, n53, n54, n58, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n71, n73, n74, n75, n76, n77, n78, n84, n85,
         n86, n87, n88, n89, n90, n91, n95, n97, n98, n99, n100, n102, n104,
         n107, n108, n109, n112, n113, n114, n115, n117, n119, n120, n121,
         n122, n123, n124, n130, n131, n132, n133, n134, n135, n136, n141,
         n143, n144, n145, n146, n147, n148, n150, n153, n154, n155, n156,
         n157, n160, n161, n163, n165, n166, n167, n168, n169, n172, n175,
         n176, n177, n178, n179, n185, n187, n188, n192, n194, n195, n197,
         n198, n199, n201, n203, n204, n205, n206, n207, n208, n214, n215,
         n216, n217, n218, n221, n225, n227, n228, n229, n230, n231, n232,
         n234, n237, n238, n239, n240, n241, n244, n245, n249, n250, n251,
         n252, n253, n254, n259, n260, n262, n271, n272, n276, n277, n278,
         n279, n280, n281, n282, n284, n286, n287, n288, n289, n293, n295,
         n296, n298, n299, n300, n304, n306, n307, n308, n309, n311, n314,
         n315, n316, n317, n319, n321, n322, n323, n324, n326, n329, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670;
  assign product[1] = a[0];

  AOI21X1 U10 ( .A(n462), .B(n670), .C(n39), .Y(n37) );
  OAI21X1 U12 ( .A(n551), .B(n662), .C(n526), .Y(n39) );
  AOI21X1 U14 ( .A(n67), .B(n638), .C(n43), .Y(n41) );
  AOI21X1 U18 ( .A(n655), .B(n58), .C(n47), .Y(n45) );
  XOR2X1 U25 ( .A(n505), .B(n541), .Y(product[29]) );
  OAI21X1 U28 ( .A(n550), .B(n664), .C(n524), .Y(n52) );
  AOI21X1 U30 ( .A(n67), .B(n642), .C(n58), .Y(n54) );
  AOI21X1 U40 ( .A(n444), .B(n457), .C(n63), .Y(n61) );
  OAI21X1 U42 ( .A(n64), .B(n663), .C(n65), .Y(n63) );
  OAI21X1 U46 ( .A(n549), .B(n563), .C(n522), .Y(n67) );
  AOI21X1 U48 ( .A(n659), .B(n84), .C(n71), .Y(n69) );
  XOR2X1 U55 ( .A(n504), .B(n540), .Y(product[27]) );
  AOI21X1 U56 ( .A(n465), .B(n670), .C(n76), .Y(n74) );
  OAI21X1 U58 ( .A(n548), .B(n662), .C(n520), .Y(n76) );
  AOI21X1 U60 ( .A(n91), .B(n643), .C(n84), .Y(n78) );
  AOI21X1 U70 ( .A(n444), .B(n461), .C(n87), .Y(n85) );
  OAI21X1 U72 ( .A(n570), .B(n663), .C(n564), .Y(n87) );
  AOI21X1 U78 ( .A(n657), .B(n104), .C(n95), .Y(n89) );
  XOR2X1 U85 ( .A(n503), .B(n539), .Y(product[25]) );
  OAI21X1 U88 ( .A(n566), .B(n664), .C(n556), .Y(n100) );
  XOR2X1 U97 ( .A(n502), .B(n538), .Y(product[24]) );
  AOI21X1 U98 ( .A(n444), .B(n108), .C(n109), .Y(n107) );
  AOI21X1 U102 ( .A(n155), .B(n482), .C(n113), .Y(n3) );
  OAI21X1 U104 ( .A(n547), .B(n561), .C(n518), .Y(n113) );
  AOI21X1 U106 ( .A(n650), .B(n130), .C(n117), .Y(n115) );
  XOR2X1 U113 ( .A(n501), .B(n537), .Y(product[23]) );
  AOI21X1 U114 ( .A(n445), .B(n460), .C(n122), .Y(n120) );
  OAI21X1 U116 ( .A(n476), .B(n157), .C(n469), .Y(n122) );
  AOI21X1 U118 ( .A(n560), .B(n641), .C(n130), .Y(n124) );
  AOI21X1 U128 ( .A(n444), .B(n459), .C(n133), .Y(n131) );
  OAI21X1 U130 ( .A(n568), .B(n157), .C(n561), .Y(n133) );
  AOI21X1 U136 ( .A(n656), .B(n150), .C(n141), .Y(n135) );
  AOI21X1 U144 ( .A(n445), .B(n458), .C(n146), .Y(n144) );
  OAI21X1 U146 ( .A(n633), .B(n157), .C(n601), .Y(n146) );
  XOR2X1 U155 ( .A(n500), .B(n536), .Y(product[20]) );
  AOI21X1 U156 ( .A(n670), .B(n559), .C(n155), .Y(n153) );
  OAI21X1 U162 ( .A(n544), .B(n585), .C(n516), .Y(n155) );
  AOI21X1 U164 ( .A(n646), .B(n172), .C(n163), .Y(n161) );
  XOR2X1 U171 ( .A(n499), .B(n535), .Y(product[19]) );
  AOI21X1 U172 ( .A(n444), .B(n528), .C(n168), .Y(n166) );
  OAI21X1 U174 ( .A(n565), .B(n585), .C(n555), .Y(n168) );
  AOI21X1 U184 ( .A(n445), .B(n176), .C(n177), .Y(n175) );
  AOI21X1 U192 ( .A(n658), .B(n192), .C(n185), .Y(n179) );
  XNOR2X1 U199 ( .A(n443), .B(n614), .Y(product[17]) );
  AOI21X1 U200 ( .A(n445), .B(n653), .C(n192), .Y(n188) );
  XOR2X1 U207 ( .A(n204), .B(n598), .Y(product[16]) );
  OAI21X1 U208 ( .A(n464), .B(n278), .C(n195), .Y(n2) );
  OAI21X1 U212 ( .A(n575), .B(n478), .C(n468), .Y(n197) );
  AOI21X1 U214 ( .A(n654), .B(n214), .C(n201), .Y(n199) );
  XOR2X1 U221 ( .A(n498), .B(n534), .Y(product[15]) );
  OAI21X1 U224 ( .A(n543), .B(n241), .C(n514), .Y(n206) );
  AOI21X1 U226 ( .A(n221), .B(n639), .C(n214), .Y(n208) );
  AOI21X1 U236 ( .A(n277), .B(n463), .C(n217), .Y(n215) );
  OAI21X1 U238 ( .A(n589), .B(n241), .C(n478), .Y(n217) );
  XOR2X1 U251 ( .A(n497), .B(n533), .Y(product[13]) );
  OAI21X1 U254 ( .A(n632), .B(n241), .C(n613), .Y(n230) );
  AOI21X1 U264 ( .A(n277), .B(n586), .C(n239), .Y(n237) );
  OAI21X1 U270 ( .A(n475), .B(n477), .C(n245), .Y(n239) );
  XOR2X1 U279 ( .A(n496), .B(n532), .Y(product[11]) );
  AOI21X1 U280 ( .A(n277), .B(n527), .C(n252), .Y(n250) );
  OAI21X1 U282 ( .A(n253), .B(n590), .C(n553), .Y(n252) );
  XOR2X1 U291 ( .A(n495), .B(n531), .Y(product[10]) );
  AOI21X1 U292 ( .A(n581), .B(n260), .C(n450), .Y(n259) );
  XNOR2X1 U307 ( .A(n581), .B(n603), .Y(product[9]) );
  AOI21X1 U308 ( .A(n277), .B(n649), .C(n276), .Y(n272) );
  XNOR2X1 U315 ( .A(n287), .B(n596), .Y(product[8]) );
  OAI21X1 U319 ( .A(n474), .B(n487), .C(n467), .Y(n280) );
  AOI21X1 U321 ( .A(n651), .B(n293), .C(n284), .Y(n282) );
  XNOR2X1 U328 ( .A(n296), .B(n604), .Y(product[7]) );
  OAI21X1 U329 ( .A(n473), .B(n314), .C(n513), .Y(n287) );
  AOI21X1 U331 ( .A(n300), .B(n640), .C(n293), .Y(n289) );
  XNOR2X1 U340 ( .A(n307), .B(n625), .Y(product[6]) );
  OAI21X1 U341 ( .A(n582), .B(n314), .C(n580), .Y(n296) );
  AOI21X1 U347 ( .A(n644), .B(n311), .C(n304), .Y(n298) );
  XOR2X1 U354 ( .A(n530), .B(n314), .Y(product[5]) );
  OAI21X1 U355 ( .A(n611), .B(n314), .C(n624), .Y(n307) );
  XNOR2X1 U364 ( .A(n322), .B(n597), .Y(product[4]) );
  OAI21X1 U366 ( .A(n635), .B(n529), .C(n511), .Y(n315) );
  AOI21X1 U368 ( .A(n326), .B(n652), .C(n319), .Y(n317) );
  OAI21X1 U376 ( .A(n610), .B(n634), .C(n622), .Y(n322) );
  INVX1 U394 ( .A(n277), .Y(n432) );
  INVX1 U395 ( .A(n277), .Y(n436) );
  OAI21X1 U396 ( .A(n432), .B(n229), .C(n433), .Y(n431) );
  INVX1 U397 ( .A(n431), .Y(n228) );
  INVX8 U398 ( .A(n230), .Y(n433) );
  INVX1 U399 ( .A(n238), .Y(n434) );
  OAI21X1 U400 ( .A(n436), .B(n205), .C(n437), .Y(n435) );
  INVX1 U401 ( .A(n435), .Y(n204) );
  INVX8 U402 ( .A(n206), .Y(n437) );
  OAI21X1 U403 ( .A(n99), .B(n442), .C(n439), .Y(n438) );
  INVX1 U404 ( .A(n438), .Y(n98) );
  INVX8 U405 ( .A(n100), .Y(n439) );
  OAI21X1 U406 ( .A(n51), .B(n442), .C(n441), .Y(n440) );
  INVX1 U407 ( .A(n440), .Y(n50) );
  INVX8 U408 ( .A(n52), .Y(n441) );
  INVX1 U409 ( .A(n445), .Y(n442) );
  INVX1 U410 ( .A(n442), .Y(n443) );
  BUFX2 U411 ( .A(n2), .Y(n444) );
  BUFX2 U412 ( .A(n2), .Y(n445) );
  AND2X2 U413 ( .A(n434), .B(n489), .Y(n194) );
  INVX1 U414 ( .A(n197), .Y(n449) );
  INVX1 U415 ( .A(n488), .Y(n448) );
  INVX1 U416 ( .A(n648), .Y(n451) );
  INVX1 U417 ( .A(n253), .Y(n446) );
  OAI21X1 U418 ( .A(n241), .B(n448), .C(n449), .Y(n447) );
  INVX1 U419 ( .A(n447), .Y(n195) );
  INVX4 U420 ( .A(n239), .Y(n241) );
  INVX1 U421 ( .A(n280), .Y(n453) );
  INVX1 U422 ( .A(n647), .Y(n455) );
  OAI21X1 U423 ( .A(n451), .B(n617), .C(n607), .Y(n450) );
  OAI21X1 U424 ( .A(n314), .B(n279), .C(n453), .Y(n452) );
  INVX1 U425 ( .A(n452), .Y(n278) );
  OAI21X1 U426 ( .A(n455), .B(n552), .C(n594), .Y(n454) );
  INVX1 U427 ( .A(n454), .Y(n245) );
  BUFX2 U428 ( .A(n2), .Y(n670) );
  AND2X2 U429 ( .A(n644), .B(n308), .Y(n456) );
  AND2X2 U430 ( .A(n509), .B(n506), .Y(n457) );
  OR2X2 U431 ( .A(n156), .B(n633), .Y(n145) );
  INVX1 U432 ( .A(n145), .Y(n458) );
  OR2X2 U433 ( .A(n156), .B(n568), .Y(n132) );
  INVX1 U434 ( .A(n132), .Y(n459) );
  OR2X2 U435 ( .A(n156), .B(n472), .Y(n121) );
  INVX1 U436 ( .A(n121), .Y(n460) );
  OR2X2 U437 ( .A(n578), .B(n570), .Y(n86) );
  INVX1 U438 ( .A(n86), .Y(n461) );
  OR2X2 U439 ( .A(n576), .B(n551), .Y(n38) );
  INVX1 U440 ( .A(n38), .Y(n462) );
  OR2X2 U441 ( .A(n240), .B(n632), .Y(n229) );
  OR2X2 U442 ( .A(n240), .B(n589), .Y(n216) );
  INVX1 U443 ( .A(n216), .Y(n463) );
  OR2X2 U444 ( .A(n240), .B(n543), .Y(n205) );
  INVX1 U445 ( .A(n194), .Y(n464) );
  OR2X2 U446 ( .A(n576), .B(n566), .Y(n99) );
  OR2X2 U447 ( .A(n577), .B(n548), .Y(n75) );
  INVX1 U448 ( .A(n75), .Y(n465) );
  OR2X2 U449 ( .A(n577), .B(n550), .Y(n51) );
  AND2X2 U450 ( .A(n638), .B(n506), .Y(n40) );
  AND2X2 U451 ( .A(a[30]), .B(a[29]), .Y(n36) );
  INVX1 U452 ( .A(n36), .Y(n466) );
  BUFX2 U453 ( .A(n282), .Y(n467) );
  BUFX2 U454 ( .A(n199), .Y(n468) );
  BUFX2 U455 ( .A(n124), .Y(n469) );
  INVX1 U456 ( .A(n281), .Y(n470) );
  INVX1 U457 ( .A(n244), .Y(n471) );
  INVX1 U458 ( .A(n123), .Y(n472) );
  OR2X2 U459 ( .A(n470), .B(n486), .Y(n279) );
  AND2X2 U460 ( .A(n640), .B(n299), .Y(n288) );
  INVX1 U461 ( .A(n288), .Y(n473) );
  AND2X2 U462 ( .A(n651), .B(n640), .Y(n281) );
  INVX1 U463 ( .A(n281), .Y(n474) );
  AND2X2 U464 ( .A(n647), .B(n587), .Y(n244) );
  INVX1 U465 ( .A(n244), .Y(n475) );
  AND2X2 U466 ( .A(n641), .B(n136), .Y(n123) );
  INVX1 U467 ( .A(n123), .Y(n476) );
  INVX1 U468 ( .A(n450), .Y(n477) );
  INVX1 U469 ( .A(n221), .Y(n478) );
  OR2X2 U470 ( .A(n557), .B(n545), .Y(n154) );
  INVX1 U471 ( .A(n154), .Y(n479) );
  INVX1 U472 ( .A(n154), .Y(n480) );
  OR2X2 U473 ( .A(n567), .B(n546), .Y(n112) );
  INVX1 U474 ( .A(n112), .Y(n481) );
  INVX1 U475 ( .A(n112), .Y(n482) );
  OR2X2 U476 ( .A(n484), .B(n471), .Y(n238) );
  INVX1 U477 ( .A(n238), .Y(n483) );
  AND2X2 U478 ( .A(n649), .B(n648), .Y(n262) );
  INVX1 U479 ( .A(n262), .Y(n484) );
  INVX1 U480 ( .A(n262), .Y(n485) );
  INVX1 U481 ( .A(n456), .Y(n486) );
  BUFX2 U482 ( .A(n298), .Y(n487) );
  OR2X2 U483 ( .A(n218), .B(n198), .Y(n542) );
  INVX1 U484 ( .A(n542), .Y(n488) );
  INVX1 U485 ( .A(n542), .Y(n489) );
  BUFX2 U486 ( .A(n250), .Y(n490) );
  BUFX2 U487 ( .A(n153), .Y(n491) );
  BUFX2 U488 ( .A(n144), .Y(n492) );
  BUFX2 U489 ( .A(n74), .Y(n493) );
  BUFX2 U490 ( .A(n37), .Y(n494) );
  BUFX2 U491 ( .A(n272), .Y(n495) );
  BUFX2 U492 ( .A(n259), .Y(n496) );
  BUFX2 U493 ( .A(n237), .Y(n497) );
  BUFX2 U494 ( .A(n215), .Y(n498) );
  BUFX2 U495 ( .A(n175), .Y(n499) );
  BUFX2 U496 ( .A(n166), .Y(n500) );
  BUFX2 U497 ( .A(n131), .Y(n501) );
  BUFX2 U498 ( .A(n120), .Y(n502) );
  BUFX2 U499 ( .A(n107), .Y(n503) );
  BUFX2 U500 ( .A(n85), .Y(n504) );
  BUFX2 U501 ( .A(n61), .Y(n505) );
  OR2X2 U502 ( .A(n569), .B(n549), .Y(n66) );
  INVX1 U503 ( .A(n66), .Y(n506) );
  INVX1 U504 ( .A(n66), .Y(n507) );
  AND2X2 U505 ( .A(a[17]), .B(a[18]), .Y(n508) );
  AND2X2 U506 ( .A(n479), .B(n481), .Y(n509) );
  OR2X2 U507 ( .A(a[24]), .B(a[23]), .Y(n510) );
  BUFX2 U508 ( .A(n317), .Y(n511) );
  INVX1 U509 ( .A(n289), .Y(n512) );
  INVX1 U510 ( .A(n512), .Y(n513) );
  BUFX2 U511 ( .A(n208), .Y(n514) );
  INVX1 U512 ( .A(n161), .Y(n515) );
  INVX1 U513 ( .A(n515), .Y(n516) );
  INVX1 U514 ( .A(n115), .Y(n517) );
  INVX1 U515 ( .A(n517), .Y(n518) );
  INVX1 U516 ( .A(n78), .Y(n519) );
  INVX1 U517 ( .A(n519), .Y(n520) );
  INVX1 U518 ( .A(n69), .Y(n521) );
  INVX1 U519 ( .A(n521), .Y(n522) );
  INVX1 U520 ( .A(n54), .Y(n523) );
  INVX1 U521 ( .A(n523), .Y(n524) );
  INVX1 U522 ( .A(n41), .Y(n525) );
  INVX1 U523 ( .A(n525), .Y(n526) );
  AND2X2 U524 ( .A(n650), .B(n641), .Y(n114) );
  OR2X2 U525 ( .A(a[23]), .B(a[22]), .Y(n650) );
  AND2X2 U526 ( .A(n659), .B(n643), .Y(n68) );
  OR2X2 U527 ( .A(a[26]), .B(a[25]), .Y(n643) );
  OR2X2 U528 ( .A(a[27]), .B(a[26]), .Y(n659) );
  OR2X2 U529 ( .A(n485), .B(n253), .Y(n251) );
  INVX1 U530 ( .A(n251), .Y(n527) );
  OR2X2 U531 ( .A(n558), .B(n565), .Y(n167) );
  INVX1 U532 ( .A(n167), .Y(n528) );
  AND2X2 U533 ( .A(n652), .B(n323), .Y(n316) );
  INVX1 U534 ( .A(n316), .Y(n529) );
  AND2X2 U535 ( .A(n624), .B(n308), .Y(n31) );
  INVX1 U536 ( .A(n31), .Y(n530) );
  AND2X2 U537 ( .A(n648), .B(n608), .Y(n26) );
  INVX1 U538 ( .A(n26), .Y(n531) );
  AND2X2 U539 ( .A(n446), .B(n553), .Y(n25) );
  INVX1 U540 ( .A(n25), .Y(n532) );
  AND2X2 U541 ( .A(n613), .B(n231), .Y(n23) );
  INVX1 U542 ( .A(n23), .Y(n533) );
  AND2X2 U543 ( .A(n628), .B(n639), .Y(n21) );
  INVX1 U544 ( .A(n21), .Y(n534) );
  AND2X2 U545 ( .A(n555), .B(n169), .Y(n17) );
  INVX1 U546 ( .A(n17), .Y(n535) );
  AND2X2 U547 ( .A(n591), .B(n646), .Y(n16) );
  INVX1 U548 ( .A(n16), .Y(n536) );
  AND2X2 U549 ( .A(n609), .B(n641), .Y(n13) );
  INVX1 U550 ( .A(n13), .Y(n537) );
  AND2X2 U551 ( .A(n618), .B(n650), .Y(n12) );
  INVX1 U552 ( .A(n12), .Y(n538) );
  AND2X2 U553 ( .A(n556), .B(n510), .Y(n11) );
  INVX1 U554 ( .A(n11), .Y(n539) );
  AND2X2 U555 ( .A(n630), .B(n643), .Y(n9) );
  INVX1 U556 ( .A(n9), .Y(n540) );
  AND2X2 U557 ( .A(n629), .B(n642), .Y(n7) );
  INVX1 U558 ( .A(n7), .Y(n541) );
  AND2X2 U559 ( .A(n639), .B(n574), .Y(n207) );
  INVX1 U560 ( .A(n207), .Y(n543) );
  AND2X2 U561 ( .A(n646), .B(n169), .Y(n160) );
  INVX1 U562 ( .A(n160), .Y(n544) );
  INVX1 U563 ( .A(n160), .Y(n545) );
  OR2X2 U564 ( .A(a[19]), .B(a[18]), .Y(n646) );
  OR2X2 U565 ( .A(a[22]), .B(a[21]), .Y(n641) );
  INVX1 U566 ( .A(n114), .Y(n546) );
  INVX1 U567 ( .A(n114), .Y(n547) );
  AND2X2 U568 ( .A(n643), .B(n90), .Y(n77) );
  INVX1 U569 ( .A(n77), .Y(n548) );
  INVX1 U570 ( .A(n68), .Y(n549) );
  AND2X2 U571 ( .A(n642), .B(n507), .Y(n53) );
  INVX1 U572 ( .A(n53), .Y(n550) );
  INVX1 U573 ( .A(n40), .Y(n551) );
  AND2X2 U574 ( .A(a[10]), .B(a[9]), .Y(n254) );
  INVX1 U575 ( .A(n254), .Y(n552) );
  INVX1 U576 ( .A(n254), .Y(n553) );
  INVX1 U577 ( .A(n508), .Y(n554) );
  INVX1 U578 ( .A(n508), .Y(n555) );
  INVX1 U579 ( .A(n102), .Y(n556) );
  AND2X2 U580 ( .A(a[23]), .B(a[24]), .Y(n102) );
  INVX1 U581 ( .A(n178), .Y(n557) );
  INVX1 U582 ( .A(n178), .Y(n558) );
  AND2X2 U583 ( .A(n658), .B(n653), .Y(n178) );
  INVX1 U584 ( .A(n156), .Y(n559) );
  INVX1 U585 ( .A(n135), .Y(n560) );
  INVX1 U586 ( .A(n560), .Y(n561) );
  INVX1 U587 ( .A(n89), .Y(n562) );
  INVX1 U588 ( .A(n562), .Y(n563) );
  INVX1 U589 ( .A(n562), .Y(n564) );
  INVX1 U590 ( .A(n169), .Y(n565) );
  OR2X2 U591 ( .A(a[18]), .B(a[17]), .Y(n169) );
  INVX1 U592 ( .A(n510), .Y(n566) );
  INVX1 U593 ( .A(n134), .Y(n567) );
  INVX1 U594 ( .A(n134), .Y(n568) );
  AND2X2 U595 ( .A(n656), .B(n147), .Y(n134) );
  INVX1 U596 ( .A(n88), .Y(n569) );
  INVX1 U597 ( .A(n88), .Y(n570) );
  AND2X2 U598 ( .A(n657), .B(n510), .Y(n88) );
  XNOR2X1 U599 ( .A(n228), .B(n571), .Y(product[14]) );
  AND2X2 U600 ( .A(n600), .B(n645), .Y(n571) );
  AOI21X1 U601 ( .A(n645), .B(n234), .C(n225), .Y(n572) );
  OR2X2 U602 ( .A(a[13]), .B(a[12]), .Y(n645) );
  AND2X2 U603 ( .A(n654), .B(n639), .Y(n573) );
  INVX1 U604 ( .A(n573), .Y(n198) );
  AND2X2 U605 ( .A(n645), .B(n231), .Y(n574) );
  INVX1 U606 ( .A(n574), .Y(n218) );
  INVX1 U607 ( .A(n573), .Y(n575) );
  INVX1 U608 ( .A(n509), .Y(n576) );
  INVX1 U609 ( .A(n509), .Y(n577) );
  INVX1 U610 ( .A(n509), .Y(n578) );
  XNOR2X1 U611 ( .A(n494), .B(n579), .Y(product[31]) );
  AND2X2 U612 ( .A(n466), .B(n660), .Y(n579) );
  INVX1 U613 ( .A(n300), .Y(n580) );
  OR2X2 U614 ( .A(a[17]), .B(a[16]), .Y(n658) );
  OR2X2 U615 ( .A(a[1]), .B(a[0]), .Y(n329) );
  OR2X2 U616 ( .A(a[10]), .B(a[11]), .Y(n647) );
  INVX1 U617 ( .A(n588), .Y(n581) );
  INVX1 U618 ( .A(n299), .Y(n582) );
  XNOR2X1 U619 ( .A(n50), .B(n583), .Y(product[30]) );
  AND2X2 U620 ( .A(n606), .B(n655), .Y(n583) );
  XNOR2X1 U621 ( .A(n490), .B(n584), .Y(product[12]) );
  AND2X2 U622 ( .A(n595), .B(n647), .Y(n584) );
  BUFX2 U623 ( .A(n179), .Y(n585) );
  INVX1 U624 ( .A(n240), .Y(n586) );
  OR2X2 U625 ( .A(a[10]), .B(a[9]), .Y(n587) );
  INVX1 U626 ( .A(n587), .Y(n253) );
  INVX1 U627 ( .A(n452), .Y(n588) );
  OR2X2 U628 ( .A(a[14]), .B(a[13]), .Y(n639) );
  INVX1 U629 ( .A(n574), .Y(n589) );
  INVX1 U630 ( .A(n450), .Y(n590) );
  XNOR2X1 U631 ( .A(n636), .B(n33), .Y(product[3]) );
  INVX2 U632 ( .A(n588), .Y(n277) );
  OR2X2 U633 ( .A(a[8]), .B(a[9]), .Y(n648) );
  AND2X2 U634 ( .A(n622), .B(n323), .Y(n33) );
  AND2X2 U635 ( .A(a[18]), .B(a[19]), .Y(n165) );
  INVX1 U636 ( .A(n165), .Y(n591) );
  AND2X2 U637 ( .A(a[20]), .B(a[21]), .Y(n143) );
  INVX1 U638 ( .A(n143), .Y(n592) );
  AND2X2 U639 ( .A(a[2]), .B(a[3]), .Y(n321) );
  INVX1 U640 ( .A(n321), .Y(n593) );
  AND2X2 U641 ( .A(a[10]), .B(a[11]), .Y(n249) );
  INVX1 U642 ( .A(n249), .Y(n594) );
  INVX1 U643 ( .A(n249), .Y(n595) );
  AND2X2 U644 ( .A(n627), .B(n651), .Y(n28) );
  INVX1 U645 ( .A(n28), .Y(n596) );
  OR2X2 U646 ( .A(a[7]), .B(a[6]), .Y(n651) );
  AND2X2 U647 ( .A(n593), .B(n652), .Y(n32) );
  INVX1 U648 ( .A(n32), .Y(n597) );
  OR2X2 U649 ( .A(a[3]), .B(a[2]), .Y(n652) );
  AND2X2 U650 ( .A(n619), .B(n654), .Y(n20) );
  INVX1 U651 ( .A(n20), .Y(n598) );
  OR2X2 U652 ( .A(a[14]), .B(a[15]), .Y(n654) );
  AND2X2 U653 ( .A(a[4]), .B(a[5]), .Y(n306) );
  INVX1 U654 ( .A(n306), .Y(n599) );
  AND2X2 U655 ( .A(a[12]), .B(a[13]), .Y(n227) );
  INVX1 U656 ( .A(n227), .Y(n600) );
  AND2X2 U657 ( .A(a[19]), .B(a[20]), .Y(n148) );
  INVX1 U658 ( .A(n148), .Y(n601) );
  BUFX2 U659 ( .A(n188), .Y(n602) );
  AND2X2 U660 ( .A(n617), .B(n649), .Y(n27) );
  INVX1 U661 ( .A(n27), .Y(n603) );
  OR2X2 U662 ( .A(a[7]), .B(a[8]), .Y(n649) );
  AND2X2 U663 ( .A(n620), .B(n640), .Y(n29) );
  INVX1 U664 ( .A(n29), .Y(n604) );
  OR2X2 U665 ( .A(a[6]), .B(a[5]), .Y(n640) );
  AND2X2 U666 ( .A(a[16]), .B(a[17]), .Y(n187) );
  INVX1 U667 ( .A(n187), .Y(n605) );
  AND2X2 U668 ( .A(a[28]), .B(a[29]), .Y(n49) );
  INVX1 U669 ( .A(n49), .Y(n606) );
  AND2X2 U670 ( .A(a[8]), .B(a[9]), .Y(n271) );
  INVX1 U671 ( .A(n271), .Y(n607) );
  INVX1 U672 ( .A(n271), .Y(n608) );
  AND2X2 U673 ( .A(a[21]), .B(a[22]), .Y(n130) );
  INVX1 U674 ( .A(n130), .Y(n609) );
  OR2X2 U675 ( .A(a[2]), .B(a[1]), .Y(n323) );
  INVX1 U676 ( .A(n323), .Y(n610) );
  OR2X2 U677 ( .A(a[4]), .B(a[3]), .Y(n308) );
  INVX1 U678 ( .A(n308), .Y(n611) );
  AND2X2 U679 ( .A(a[11]), .B(a[12]), .Y(n232) );
  INVX1 U680 ( .A(n232), .Y(n612) );
  INVX1 U681 ( .A(n232), .Y(n613) );
  AND2X2 U682 ( .A(n631), .B(n653), .Y(n19) );
  INVX1 U683 ( .A(n19), .Y(n614) );
  OR2X2 U684 ( .A(a[16]), .B(a[15]), .Y(n653) );
  AND2X2 U685 ( .A(a[26]), .B(a[27]), .Y(n73) );
  INVX1 U686 ( .A(n73), .Y(n615) );
  AND2X2 U687 ( .A(a[24]), .B(a[25]), .Y(n97) );
  INVX1 U688 ( .A(n97), .Y(n616) );
  AND2X2 U689 ( .A(a[7]), .B(a[8]), .Y(n276) );
  INVX1 U690 ( .A(n276), .Y(n617) );
  AND2X2 U691 ( .A(a[22]), .B(a[23]), .Y(n119) );
  INVX1 U692 ( .A(n119), .Y(n618) );
  AND2X2 U693 ( .A(a[14]), .B(a[15]), .Y(n203) );
  INVX1 U694 ( .A(n203), .Y(n619) );
  AND2X2 U695 ( .A(a[5]), .B(a[6]), .Y(n295) );
  INVX1 U696 ( .A(n295), .Y(n620) );
  AND2X2 U697 ( .A(a[2]), .B(a[1]), .Y(n324) );
  INVX1 U698 ( .A(n324), .Y(n621) );
  INVX1 U699 ( .A(n324), .Y(n622) );
  AND2X2 U700 ( .A(a[4]), .B(a[3]), .Y(n309) );
  INVX1 U701 ( .A(n309), .Y(n623) );
  INVX1 U702 ( .A(n309), .Y(n624) );
  AND2X2 U703 ( .A(n599), .B(n644), .Y(n30) );
  INVX1 U704 ( .A(n30), .Y(n625) );
  AND2X2 U705 ( .A(a[7]), .B(a[6]), .Y(n286) );
  INVX1 U706 ( .A(n286), .Y(n626) );
  INVX1 U707 ( .A(n286), .Y(n627) );
  AND2X2 U708 ( .A(a[13]), .B(a[14]), .Y(n214) );
  INVX1 U709 ( .A(n214), .Y(n628) );
  AND2X2 U710 ( .A(a[27]), .B(a[28]), .Y(n60) );
  INVX1 U711 ( .A(n60), .Y(n629) );
  AND2X2 U712 ( .A(a[25]), .B(a[26]), .Y(n84) );
  INVX1 U713 ( .A(n84), .Y(n630) );
  AND2X2 U714 ( .A(a[15]), .B(a[16]), .Y(n192) );
  INVX1 U715 ( .A(n192), .Y(n631) );
  OR2X2 U716 ( .A(a[12]), .B(a[11]), .Y(n231) );
  INVX1 U717 ( .A(n231), .Y(n632) );
  OR2X2 U718 ( .A(a[20]), .B(a[19]), .Y(n147) );
  INVX1 U719 ( .A(n147), .Y(n633) );
  AND2X2 U720 ( .A(a[1]), .B(a[0]), .Y(n1) );
  INVX1 U721 ( .A(n1), .Y(n634) );
  INVX1 U722 ( .A(n1), .Y(n635) );
  INVX1 U723 ( .A(n1), .Y(n636) );
  AND2X2 U724 ( .A(n634), .B(n329), .Y(product[2]) );
  OR2X2 U725 ( .A(a[4]), .B(a[5]), .Y(n644) );
  INVX1 U726 ( .A(n578), .Y(n108) );
  INVX1 U727 ( .A(n480), .Y(n156) );
  INVX1 U728 ( .A(n483), .Y(n240) );
  INVX1 U729 ( .A(n507), .Y(n64) );
  INVX1 U730 ( .A(n485), .Y(n260) );
  INVX1 U731 ( .A(n155), .Y(n157) );
  INVX1 U732 ( .A(n67), .Y(n65) );
  INVX1 U733 ( .A(n585), .Y(n177) );
  INVX1 U734 ( .A(n615), .Y(n71) );
  INVX1 U735 ( .A(n591), .Y(n163) );
  INVX1 U736 ( .A(n554), .Y(n172) );
  INVX1 U737 ( .A(n605), .Y(n185) );
  INVX1 U738 ( .A(n600), .Y(n225) );
  INVX1 U739 ( .A(n612), .Y(n234) );
  INVX1 U740 ( .A(n592), .Y(n141) );
  INVX1 U741 ( .A(n601), .Y(n150) );
  INVX1 U742 ( .A(n616), .Y(n95) );
  INVX1 U743 ( .A(n556), .Y(n104) );
  INVX1 U744 ( .A(n593), .Y(n319) );
  INVX1 U745 ( .A(n568), .Y(n136) );
  INVX1 U746 ( .A(n569), .Y(n90) );
  INVX1 U747 ( .A(n599), .Y(n304) );
  INVX1 U748 ( .A(n623), .Y(n311) );
  INVX1 U749 ( .A(n663), .Y(n109) );
  INVX1 U750 ( .A(n558), .Y(n176) );
  INVX1 U751 ( .A(n45), .Y(n43) );
  INVX1 U752 ( .A(n619), .Y(n201) );
  INVX1 U753 ( .A(n572), .Y(n221) );
  INVX1 U754 ( .A(n564), .Y(n91) );
  INVX1 U755 ( .A(n621), .Y(n326) );
  INVX1 U756 ( .A(n620), .Y(n293) );
  INVX1 U757 ( .A(n629), .Y(n58) );
  INVX1 U758 ( .A(n618), .Y(n117) );
  INVX1 U759 ( .A(n626), .Y(n284) );
  INVX1 U760 ( .A(n606), .Y(n47) );
  AND2X1 U761 ( .A(n655), .B(n642), .Y(n638) );
  OR2X1 U762 ( .A(a[28]), .B(a[27]), .Y(n642) );
  OR2X1 U763 ( .A(a[29]), .B(a[28]), .Y(n655) );
  OR2X1 U764 ( .A(a[21]), .B(a[20]), .Y(n656) );
  OR2X1 U765 ( .A(a[25]), .B(a[24]), .Y(n657) );
  OR2X1 U766 ( .A(a[29]), .B(a[30]), .Y(n660) );
  INVX1 U767 ( .A(n487), .Y(n300) );
  INVX1 U768 ( .A(n315), .Y(n314) );
  INVX1 U769 ( .A(n486), .Y(n299) );
  INVX1 U770 ( .A(n3), .Y(n661) );
  INVX1 U771 ( .A(n661), .Y(n662) );
  INVX1 U772 ( .A(n661), .Y(n663) );
  INVX1 U773 ( .A(n661), .Y(n664) );
  XNOR2X1 U774 ( .A(n493), .B(n665), .Y(product[28]) );
  AND2X2 U775 ( .A(n615), .B(n659), .Y(n665) );
  XNOR2X1 U776 ( .A(n98), .B(n666), .Y(product[26]) );
  AND2X2 U777 ( .A(n616), .B(n657), .Y(n666) );
  XNOR2X1 U778 ( .A(n491), .B(n667), .Y(product[21]) );
  AND2X2 U779 ( .A(n601), .B(n147), .Y(n667) );
  XNOR2X1 U780 ( .A(n492), .B(n668), .Y(product[22]) );
  AND2X2 U781 ( .A(n592), .B(n656), .Y(n668) );
  XNOR2X1 U782 ( .A(n602), .B(n669), .Y(product[18]) );
  AND2X2 U783 ( .A(n605), .B(n658), .Y(n669) );
endmodule


module maze_router_DW01_add_10 ( A, B, CI, SUM, CO );
  input [179:0] A;
  input [179:0] B;
  output [179:0] SUM;
  input CI;
  output CO;
  wire   n7, n15, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30,
         n32, n33, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n48,
         n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n146, n147, n148, n149, n150,
         n151, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n172, n173, n174, n176,
         n177, n178, n180, n181, n182, n183, n184, n185, n186, n188, n191,
         n194, n195, n196, n199, n200, n202, n204, n205, n206, n207, n208,
         n210, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n228, n229, n230, n231, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n252, n253, n254, n255, n257, n258, n259, n260,
         n261, n262, n265, n267, n268, n269, n270, n271, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n285, n288, n289, n290,
         n291, n292, n293, n294, n295, n298, n299, n300, n301, n302, n303,
         n304, n305, n307, n309, n310, n311, n312, n313, n314, n315, n318,
         n319, n320, n321, n322, n323, n324, n325, n327, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n343, n344, n345, n346,
         n347, n348, n349, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n376, n377, n378, n379, n380, n381, n382, n383, n386, n387, n388,
         n389, n390, n391, n392, n395, n396, n397, n398, n399, n400, n401,
         n404, n405, n406, n407, n408, n409, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n441, n443,
         n444, n445, n446, n450, n451, n453, n454, n455, n456, n457, n458,
         n459, n461, n464, n465, n466, n467, n468, n469, n470, n471, n474,
         n475, n476, n477, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n552, n553, n554,
         n555, n556, n557, n558, n562, n563, n564, n565, n566, n567, n568,
         n571, n572, n573, n574, n575, n576, n577, n580, n581, n584, n585,
         n587, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n604, n605, n606, n607, n608, n609, n610, n613, n614, n615,
         n616, n617, n618, n622, n623, n624, n625, n626, n627, n630, n633,
         n634, n635, n636, n637, n638, n639, n640, n644, n645, n646, n647,
         n648, n649, n650, n653, n654, n655, n656, n657, n658, n662, n663,
         n668, n669, n670, n671, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n687, n688, n689, n690, n691, n692, n695, n697, n698,
         n699, n700, n705, n708, n709, n711, n714, n715, n716, n717, n718,
         n719, n720, n725, n726, n727, n728, n729, n732, n733, n734, n736,
         n737, n738, n740, n741, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n856, n857, n858, n859, n860, n861, n862, n863, n865, n868, n869,
         n870, n871, n873, n874, n875, n876, n877, n878, n879, n880, n884,
         n885, n887, n888, n889, n890, n891, n892, n893, n894, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n910, n911, n912,
         n913, n914, n915, n918, n919, n921, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n938, n939, n940, n941, n942,
         n943, n944, n945, n947, n950, n951, n952, n953, n954, n955, n956,
         n959, n961, n962, n963, n964, n965, n967, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n984, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n999,
         n1001, n1002, n1003, n1004, n1005, n1006, n1009, n1010, n1011, n1012,
         n1013, n1014, n1016, n1017, n1018, n1019, n1020, n1021, n1024, n1025,
         n1027, n1028, n1029, n1030, n1031, n1032, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1059, n1060, n1061, n1064, n1065,
         n1067, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1082, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1095, n1097, n1098, n1099, n1100, n1101, n1102,
         n1107, n1108, n1109, n1112, n1113, n1114, n1115, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1130, n1131, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1145, n1146, n1147, n1148, n1149,
         n1153, n1155, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1177, n1178, n1179, n1180, n1182,
         n1183, n1184, n1185, n1186, n1189, n1191, n1192, n1193, n1194, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1267, n1268, n1269, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1286,
         n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1319, n1320, n1321, n1322, n1323, n1324, n1328, n1329,
         n1332, n1333, n1335, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1361, n1363, n1364, n1365, n1366, n1370, n1371, n1372, n1373,
         n1375, n1378, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1393, n1394, n1395, n1396, n1397, n1398, n1401, n1403, n1404,
         n1405, n1406, n1411, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1435, n1436, n1437, n1438, n1439, n1440, n1443, n1444,
         n1445, n1446, n1447, n1448, n1453, n1456, n1457, n1459, n1462, n1463,
         n1465, n1466, n1467, n1468, n1469, n1473, n1474, n1475, n1476, n1477,
         n1481, n1482, n1484, n1485, n1486, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1505, n1506, n1507, n1508, n1509, n1510, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1564, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1624, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1635, n1636, n1637, n1638, n1641, n1642, n1643, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1670, n1671, n1672, n1673,
         n1676, n1678, n1679, n1680, n1681, n1682, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1697, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1710, n1712, n1713, n1714,
         n1715, n1717, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1752, n1753, n1754, n1755, n1758, n1760, n1764, n1765, n1769, n1770,
         n1772, n1773, n1774, n1775, n1776, n1777, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1797, n1798, n1799, n1800, n1803, n1804, n1805,
         n1806, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1832, n1833, n1834, n1835,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1890, n1891, n1893, n1894, n1895, n1896, n1897, n1898,
         n1900, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1915,
         n1916, n1917, n1918, n1919, n1922, n1923, n1924, n1925, n1926, n1927,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1942,
         n1943, n1945, n1947, n1948, n1951, n1953, n1954, n1955, n1956, n1961,
         n1964, n1965, n1966, n1967, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1980, n1982, n1983, n1985, n1989, n1990, n1993, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2009, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2023, n2024, n2025, n2026, n2027, n2030, n2032, n2033, n2034, n2035,
         n2036, n2040, n2041, n2042, n2043, n2044, n2045, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2071, n2072, n2074, n2075, n2078, n2079,
         n2080, n2081, n2082, n2083, n2087, n2088, n2091, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2101, n2102, n2103, n2105, n2107, n2111,
         n2113, n2114, n2115, n2117, n2118, n2119, n2120, n2121, n2123, n2125,
         n2126, n2127, n2128, n2129, n2130, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2143, n2144, n2148, n2149, n2151, n2152,
         n2155, n2156, n2158, n2160, n2164, n2166, n2167, n2173, n2176, n2180,
         n2181, n2182, n2184, n2187, n2188, n2189, n2191, n2195, n2199, n2200,
         n2202, n2203, n2204, n2205, n2207, n2208, n2211, n2214, n2216, n2218,
         n2221, n2222, n2224, n2225, n2226, n2227, n2228, n2229, n2231, n2232,
         n2233, n2236, n2240, n2242, n2244, n2248, n2250, n2251, n2253, n2258,
         n2260, n2264, n2266, n2268, n2269, n2270, n2275, n2282, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794;

  XOR2X1 U18 ( .A(n3720), .B(n4132), .Y(SUM[179]) );
  XOR2X1 U23 ( .A(n3719), .B(n4131), .Y(SUM[178]) );
  AOI21X1 U24 ( .A(n2888), .B(n4782), .C(n202), .Y(n200) );
  AOI21X1 U28 ( .A(n4741), .B(n2949), .C(n206), .Y(n204) );
  OAI21X1 U30 ( .A(n3231), .B(n4313), .C(n3865), .Y(n206) );
  AOI21X1 U32 ( .A(n219), .B(n4783), .C(n210), .Y(n208) );
  XOR2X1 U39 ( .A(n3718), .B(n4130), .Y(SUM[177]) );
  AOI21X1 U40 ( .A(n4791), .B(n3144), .C(n215), .Y(n213) );
  OAI21X1 U42 ( .A(n216), .B(n3554), .C(n217), .Y(n215) );
  OAI21X1 U46 ( .A(n3492), .B(n4530), .C(n3143), .Y(n219) );
  XOR2X1 U51 ( .A(n3717), .B(n4129), .Y(SUM[176]) );
  AOI21X1 U52 ( .A(n2889), .B(n3142), .C(n224), .Y(n222) );
  OAI21X1 U54 ( .A(n4633), .B(n3554), .C(n3493), .Y(n224) );
  XOR2X1 U61 ( .A(n3716), .B(n4128), .Y(SUM[175]) );
  AOI21X1 U62 ( .A(n2863), .B(n230), .C(n231), .Y(n229) );
  AOI21X1 U66 ( .A(n4790), .B(n234), .C(n235), .Y(n233) );
  AOI21X1 U70 ( .A(n325), .B(n3572), .C(n239), .Y(n237) );
  OAI21X1 U72 ( .A(n3602), .B(n4343), .C(n3864), .Y(n239) );
  AOI21X1 U74 ( .A(n265), .B(n3561), .C(n243), .Y(n241) );
  OAI21X1 U76 ( .A(n4219), .B(n4529), .C(n3140), .Y(n243) );
  XOR2X1 U81 ( .A(n3715), .B(n4127), .Y(SUM[174]) );
  AOI21X1 U82 ( .A(n4791), .B(n3139), .C(n248), .Y(n246) );
  OAI21X1 U84 ( .A(n4632), .B(n3553), .C(n4577), .Y(n248) );
  XOR2X1 U91 ( .A(n3714), .B(n4126), .Y(SUM[173]) );
  AOI21X1 U92 ( .A(n2888), .B(n254), .C(n255), .Y(n253) );
  AOI21X1 U96 ( .A(n4740), .B(n4288), .C(n259), .Y(n257) );
  OAI21X1 U98 ( .A(n3394), .B(n327), .C(n3862), .Y(n259) );
  AOI21X1 U100 ( .A(n285), .B(n4549), .C(n265), .Y(n261) );
  OAI21X1 U104 ( .A(n3218), .B(n3524), .C(n3365), .Y(n265) );
  XOR2X1 U109 ( .A(n3713), .B(n4125), .Y(SUM[172]) );
  AOI21X1 U110 ( .A(n4791), .B(n3137), .C(n270), .Y(n268) );
  OAI21X1 U112 ( .A(n4630), .B(n3552), .C(n3523), .Y(n270) );
  XOR2X1 U119 ( .A(n3712), .B(n4124), .Y(SUM[171]) );
  AOI21X1 U120 ( .A(n2888), .B(n276), .C(n277), .Y(n275) );
  AOI21X1 U124 ( .A(n4741), .B(n4287), .C(n281), .Y(n279) );
  OAI21X1 U126 ( .A(n4628), .B(n327), .C(n4343), .Y(n281) );
  AOI21X1 U132 ( .A(n309), .B(n3564), .C(n289), .Y(n283) );
  OAI21X1 U134 ( .A(n4218), .B(n4528), .C(n3136), .Y(n289) );
  XOR2X1 U139 ( .A(n3711), .B(n4123), .Y(SUM[170]) );
  AOI21X1 U140 ( .A(n2864), .B(n3135), .C(n294), .Y(n292) );
  OAI21X1 U142 ( .A(n4626), .B(n3551), .C(n4576), .Y(n294) );
  XOR2X1 U149 ( .A(n3710), .B(n4122), .Y(SUM[169]) );
  AOI21X1 U150 ( .A(n2864), .B(n300), .C(n301), .Y(n299) );
  AOI21X1 U154 ( .A(n4790), .B(n2948), .C(n305), .Y(n303) );
  OAI21X1 U156 ( .A(n3753), .B(n327), .C(n307), .Y(n305) );
  OAI21X1 U160 ( .A(n3490), .B(n4527), .C(n3134), .Y(n309) );
  AOI21X1 U166 ( .A(n4791), .B(n3133), .C(n314), .Y(n312) );
  OAI21X1 U168 ( .A(n4624), .B(n3550), .C(n3491), .Y(n314) );
  XOR2X1 U175 ( .A(n3709), .B(n4121), .Y(SUM[167]) );
  AOI21X1 U176 ( .A(n4791), .B(n320), .C(n321), .Y(n319) );
  AOI21X1 U180 ( .A(n4741), .B(n4599), .C(n325), .Y(n323) );
  OAI21X1 U186 ( .A(n3356), .B(n3547), .C(n3861), .Y(n325) );
  AOI21X1 U188 ( .A(n353), .B(n3260), .C(n333), .Y(n331) );
  OAI21X1 U190 ( .A(n2918), .B(n4525), .C(n3131), .Y(n333) );
  AOI21X1 U196 ( .A(n2888), .B(n3130), .C(n338), .Y(n336) );
  OAI21X1 U198 ( .A(n4622), .B(n3549), .C(n2918), .Y(n338) );
  XOR2X1 U205 ( .A(n3708), .B(n4120), .Y(SUM[165]) );
  AOI21X1 U206 ( .A(n2888), .B(n344), .C(n345), .Y(n343) );
  AOI21X1 U210 ( .A(n4741), .B(n2947), .C(n349), .Y(n347) );
  OAI21X1 U212 ( .A(n352), .B(n4586), .C(n351), .Y(n349) );
  OAI21X1 U216 ( .A(n3217), .B(n4523), .C(n3129), .Y(n353) );
  XOR2X1 U221 ( .A(n3707), .B(n4119), .Y(SUM[164]) );
  AOI21X1 U222 ( .A(n2876), .B(n3128), .C(n358), .Y(n356) );
  OAI21X1 U224 ( .A(n4619), .B(n3548), .C(n3217), .Y(n358) );
  AOI21X1 U232 ( .A(n2888), .B(n364), .C(n365), .Y(n363) );
  AOI21X1 U236 ( .A(n4740), .B(n368), .C(n369), .Y(n367) );
  AOI21X1 U244 ( .A(n395), .B(n3570), .C(n377), .Y(n371) );
  OAI21X1 U246 ( .A(n3488), .B(n4522), .C(n3126), .Y(n377) );
  XOR2X1 U251 ( .A(n3706), .B(n4118), .Y(SUM[162]) );
  AOI21X1 U252 ( .A(n2868), .B(n3125), .C(n382), .Y(n380) );
  OAI21X1 U254 ( .A(n4618), .B(n3546), .C(n3489), .Y(n382) );
  XOR2X1 U261 ( .A(n3705), .B(n4117), .Y(SUM[161]) );
  AOI21X1 U262 ( .A(n4791), .B(n388), .C(n389), .Y(n387) );
  AOI21X1 U266 ( .A(n4790), .B(n4547), .C(n395), .Y(n391) );
  OAI21X1 U270 ( .A(n4574), .B(n4520), .C(n4209), .Y(n395) );
  XOR2X1 U275 ( .A(n3704), .B(n4116), .Y(SUM[160]) );
  AOI21X1 U276 ( .A(n2888), .B(n2946), .C(n400), .Y(n398) );
  OAI21X1 U278 ( .A(n4616), .B(n409), .C(n4575), .Y(n400) );
  XOR2X1 U285 ( .A(n3703), .B(n4115), .Y(SUM[159]) );
  AOI21X1 U286 ( .A(n4791), .B(n406), .C(n4740), .Y(n405) );
  OAI21X1 U292 ( .A(n3123), .B(n3540), .C(n3168), .Y(n407) );
  AOI21X1 U294 ( .A(n501), .B(n2945), .C(n415), .Y(n413) );
  OAI21X1 U296 ( .A(n3600), .B(n3543), .C(n3859), .Y(n415) );
  AOI21X1 U298 ( .A(n441), .B(n3258), .C(n419), .Y(n417) );
  OAI21X1 U300 ( .A(n4572), .B(n4519), .C(n3122), .Y(n419) );
  XOR2X1 U305 ( .A(n3702), .B(n4114), .Y(SUM[158]) );
  AOI21X1 U306 ( .A(n2889), .B(n3949), .C(n424), .Y(n422) );
  OAI21X1 U308 ( .A(n4614), .B(n3545), .C(n4573), .Y(n424) );
  XOR2X1 U315 ( .A(n3701), .B(n4113), .Y(SUM[157]) );
  AOI21X1 U316 ( .A(n2864), .B(n430), .C(n431), .Y(n429) );
  AOI21X1 U320 ( .A(n4684), .B(n3121), .C(n435), .Y(n433) );
  OAI21X1 U322 ( .A(n4312), .B(n503), .C(n3857), .Y(n435) );
  AOI21X1 U324 ( .A(n461), .B(n4545), .C(n441), .Y(n437) );
  OAI21X1 U328 ( .A(n3976), .B(n4570), .C(n3119), .Y(n441) );
  XOR2X1 U333 ( .A(n3700), .B(n4112), .Y(SUM[156]) );
  AOI21X1 U334 ( .A(n2869), .B(n2944), .C(n446), .Y(n444) );
  OAI21X1 U336 ( .A(n4365), .B(n3544), .C(n4571), .Y(n446) );
  AOI21X1 U344 ( .A(n2888), .B(n454), .C(n453), .Y(n451) );
  AOI21X1 U348 ( .A(n4682), .B(n4273), .C(n457), .Y(n455) );
  OAI21X1 U350 ( .A(n4401), .B(n503), .C(n4342), .Y(n457) );
  AOI21X1 U356 ( .A(n485), .B(n3890), .C(n465), .Y(n459) );
  OAI21X1 U358 ( .A(n4568), .B(n4517), .C(n4165), .Y(n465) );
  XOR2X1 U363 ( .A(n3699), .B(n4111), .Y(SUM[154]) );
  AOI21X1 U364 ( .A(n4791), .B(n3948), .C(n470), .Y(n468) );
  OAI21X1 U366 ( .A(n4612), .B(n3542), .C(n4569), .Y(n470) );
  XOR2X1 U373 ( .A(n3698), .B(n4110), .Y(SUM[153]) );
  AOI21X1 U374 ( .A(n2888), .B(n476), .C(n477), .Y(n475) );
  AOI21X1 U378 ( .A(n4682), .B(n3116), .C(n481), .Y(n479) );
  OAI21X1 U380 ( .A(n482), .B(n503), .C(n483), .Y(n481) );
  OAI21X1 U384 ( .A(n4566), .B(n4515), .C(n3114), .Y(n485) );
  XOR2X1 U389 ( .A(n3697), .B(n4109), .Y(SUM[152]) );
  AOI21X1 U390 ( .A(n4738), .B(n3947), .C(n490), .Y(n488) );
  OAI21X1 U392 ( .A(n4241), .B(n4610), .C(n4567), .Y(n490) );
  XOR2X1 U399 ( .A(n3696), .B(n4108), .Y(SUM[151]) );
  AOI21X1 U400 ( .A(n2889), .B(n496), .C(n497), .Y(n495) );
  AOI21X1 U404 ( .A(n4683), .B(n4597), .C(n501), .Y(n499) );
  OAI21X1 U410 ( .A(n4311), .B(n3541), .C(n3856), .Y(n501) );
  AOI21X1 U412 ( .A(n529), .B(n3322), .C(n509), .Y(n507) );
  OAI21X1 U414 ( .A(n3112), .B(n4513), .C(n4208), .Y(n509) );
  AOI21X1 U420 ( .A(n2888), .B(n3946), .C(n514), .Y(n512) );
  OAI21X1 U422 ( .A(n4240), .B(n4369), .C(n3112), .Y(n514) );
  XOR2X1 U429 ( .A(n3695), .B(n4107), .Y(SUM[149]) );
  AOI21X1 U430 ( .A(n2888), .B(n520), .C(n521), .Y(n519) );
  AOI21X1 U434 ( .A(n4683), .B(n2943), .C(n525), .Y(n523) );
  OAI21X1 U436 ( .A(n526), .B(n4585), .C(n527), .Y(n525) );
  OAI21X1 U440 ( .A(n4362), .B(n4511), .C(n4207), .Y(n529) );
  AOI21X1 U446 ( .A(n4791), .B(n3945), .C(n534), .Y(n532) );
  OAI21X1 U448 ( .A(n4239), .B(n4608), .C(n4363), .Y(n534) );
  XOR2X1 U455 ( .A(n3694), .B(n4106), .Y(SUM[147]) );
  AOI21X1 U456 ( .A(n4791), .B(n540), .C(n541), .Y(n539) );
  AOI21X1 U460 ( .A(n4684), .B(n544), .C(n545), .Y(n543) );
  AOI21X1 U468 ( .A(n571), .B(n3256), .C(n553), .Y(n547) );
  OAI21X1 U470 ( .A(n2942), .B(n4509), .C(n4206), .Y(n553) );
  XOR2X1 U475 ( .A(n3693), .B(n4105), .Y(SUM[146]) );
  AOI21X1 U476 ( .A(n2888), .B(n3944), .C(n558), .Y(n556) );
  OAI21X1 U478 ( .A(n4238), .B(n4371), .C(n2942), .Y(n558) );
  XOR2X1 U485 ( .A(n3692), .B(n4104), .Y(SUM[145]) );
  AOI21X1 U486 ( .A(n2868), .B(n564), .C(n565), .Y(n563) );
  AOI21X1 U490 ( .A(n4684), .B(n4544), .C(n571), .Y(n567) );
  OAI21X1 U494 ( .A(n4507), .B(n4564), .C(n4205), .Y(n571) );
  XOR2X1 U499 ( .A(n3691), .B(n4103), .Y(SUM[144]) );
  AOI21X1 U500 ( .A(n2869), .B(n3943), .C(n576), .Y(n574) );
  OAI21X1 U502 ( .A(n4584), .B(n4605), .C(n4565), .Y(n576) );
  XOR2X1 U509 ( .A(n3690), .B(n4102), .Y(SUM[143]) );
  AOI21X1 U510 ( .A(n2888), .B(n584), .C(n4683), .Y(n581) );
  AOI21X1 U518 ( .A(n669), .B(n3110), .C(n591), .Y(n585) );
  OAI21X1 U520 ( .A(n3109), .B(n3506), .C(n3854), .Y(n591) );
  AOI21X1 U522 ( .A(n613), .B(n3108), .C(n595), .Y(n593) );
  OAI21X1 U524 ( .A(n3486), .B(n3107), .C(n3106), .Y(n595) );
  AOI21X1 U530 ( .A(n4791), .B(n3942), .C(n600), .Y(n598) );
  OAI21X1 U532 ( .A(n4374), .B(n3539), .C(n3487), .Y(n600) );
  XOR2X1 U539 ( .A(n3689), .B(n4101), .Y(SUM[141]) );
  AOI21X1 U540 ( .A(n2888), .B(n606), .C(n607), .Y(n605) );
  AOI21X1 U544 ( .A(n625), .B(n4543), .C(n613), .Y(n609) );
  OAI21X1 U548 ( .A(n3484), .B(n2882), .C(n3104), .Y(n613) );
  XOR2X1 U553 ( .A(n3688), .B(n4100), .Y(SUM[140]) );
  AOI21X1 U554 ( .A(n2869), .B(n3941), .C(n618), .Y(n616) );
  OAI21X1 U556 ( .A(n4385), .B(n627), .C(n3485), .Y(n618) );
  XOR2X1 U563 ( .A(n3687), .B(n4099), .Y(SUM[139]) );
  AOI21X1 U564 ( .A(n4738), .B(n4330), .C(n625), .Y(n623) );
  OAI21X1 U570 ( .A(n4588), .B(n671), .C(n4290), .Y(n625) );
  AOI21X1 U574 ( .A(n653), .B(n3102), .C(n635), .Y(n633) );
  OAI21X1 U576 ( .A(n3482), .B(n3101), .C(n3100), .Y(n635) );
  XOR2X1 U581 ( .A(n3686), .B(n4098), .Y(SUM[138]) );
  AOI21X1 U582 ( .A(n2888), .B(n3940), .C(n640), .Y(n638) );
  OAI21X1 U584 ( .A(n4415), .B(n3538), .C(n4563), .Y(n640) );
  XOR2X1 U591 ( .A(n3685), .B(n4097), .Y(SUM[137]) );
  AOI21X1 U592 ( .A(n2888), .B(n646), .C(n647), .Y(n645) );
  AOI21X1 U596 ( .A(n4744), .B(n4542), .C(n653), .Y(n649) );
  OAI21X1 U600 ( .A(n4466), .B(n3522), .C(n3099), .Y(n653) );
  XOR2X1 U605 ( .A(n3684), .B(n4096), .Y(SUM[136]) );
  AOI21X1 U606 ( .A(n4791), .B(n3939), .C(n658), .Y(n656) );
  OAI21X1 U608 ( .A(n4393), .B(n671), .C(n4562), .Y(n658) );
  XOR2X1 U615 ( .A(n3683), .B(n4095), .Y(SUM[135]) );
  AOI21X1 U616 ( .A(n2876), .B(n4589), .C(n4744), .Y(n663) );
  OAI21X1 U626 ( .A(n3598), .B(n3537), .C(n3852), .Y(n669) );
  AOI21X1 U628 ( .A(n695), .B(n3098), .C(n677), .Y(n675) );
  OAI21X1 U630 ( .A(n2923), .B(n4465), .C(n3096), .Y(n677) );
  XOR2X1 U635 ( .A(n3682), .B(n4094), .Y(SUM[134]) );
  AOI21X1 U636 ( .A(n2863), .B(n3938), .C(n682), .Y(n680) );
  OAI21X1 U638 ( .A(n4237), .B(n4396), .C(n2923), .Y(n682) );
  XOR2X1 U645 ( .A(n3681), .B(n4093), .Y(SUM[133]) );
  AOI21X1 U646 ( .A(n2876), .B(n688), .C(n689), .Y(n687) );
  AOI21X1 U650 ( .A(n711), .B(n4540), .C(n695), .Y(n691) );
  OAI21X1 U654 ( .A(n2917), .B(n4506), .C(n3095), .Y(n695) );
  XOR2X1 U659 ( .A(n3680), .B(n4092), .Y(SUM[132]) );
  AOI21X1 U660 ( .A(n4738), .B(n3937), .C(n700), .Y(n698) );
  OAI21X1 U662 ( .A(n4583), .B(n4469), .C(n2917), .Y(n700) );
  XOR2X1 U669 ( .A(n3679), .B(n4091), .Y(SUM[131]) );
  AOI21X1 U670 ( .A(n4791), .B(n708), .C(n711), .Y(n705) );
  AOI21X1 U678 ( .A(n727), .B(n3319), .C(n715), .Y(n709) );
  OAI21X1 U680 ( .A(n3470), .B(n3094), .C(n3093), .Y(n715) );
  XOR2X1 U685 ( .A(n3678), .B(n4090), .Y(SUM[130]) );
  AOI21X1 U686 ( .A(n4791), .B(n3936), .C(n720), .Y(n718) );
  OAI21X1 U688 ( .A(n4419), .B(n729), .C(n3471), .Y(n720) );
  XOR2X1 U695 ( .A(n3677), .B(n4089), .Y(SUM[129]) );
  AOI21X1 U696 ( .A(n4791), .B(n4329), .C(n4672), .Y(n725) );
  OAI21X1 U702 ( .A(n4353), .B(n4504), .C(n4204), .Y(n727) );
  XNOR2X1 U707 ( .A(n4691), .B(n4015), .Y(SUM[128]) );
  AOI21X1 U708 ( .A(n2863), .B(n737), .C(n736), .Y(n734) );
  XOR2X1 U715 ( .A(n3676), .B(n4088), .Y(SUM[127]) );
  OAI21X1 U716 ( .A(n3216), .B(n2853), .C(n3167), .Y(n15) );
  AOI21X1 U718 ( .A(n2899), .B(n2904), .C(n743), .Y(n741) );
  OAI21X1 U720 ( .A(n3739), .B(n3462), .C(n3850), .Y(n743) );
  AOI21X1 U722 ( .A(n863), .B(n3092), .C(n747), .Y(n745) );
  OAI21X1 U724 ( .A(n3403), .B(n4340), .C(n3848), .Y(n747) );
  AOI21X1 U726 ( .A(n779), .B(n4286), .C(n751), .Y(n749) );
  OAI21X1 U728 ( .A(n4463), .B(n3520), .C(n3090), .Y(n751) );
  XOR2X1 U733 ( .A(n3675), .B(n4087), .Y(SUM[126]) );
  AOI21X1 U734 ( .A(n4776), .B(n3089), .C(n756), .Y(n754) );
  OAI21X1 U736 ( .A(n3460), .B(n4793), .C(n3166), .Y(n756) );
  AOI21X1 U738 ( .A(n4718), .B(n4272), .C(n760), .Y(n758) );
  OAI21X1 U740 ( .A(n4310), .B(n865), .C(n3847), .Y(n760) );
  AOI21X1 U742 ( .A(n809), .B(n4256), .C(n764), .Y(n762) );
  OAI21X1 U744 ( .A(n4382), .B(n781), .C(n4561), .Y(n764) );
  XOR2X1 U751 ( .A(n3674), .B(n4086), .Y(SUM[125]) );
  AOI21X1 U752 ( .A(n4659), .B(n3088), .C(n771), .Y(n769) );
  OAI21X1 U754 ( .A(n3458), .B(n2845), .C(n3165), .Y(n771) );
  AOI21X1 U756 ( .A(n4718), .B(n4270), .C(n775), .Y(n773) );
  OAI21X1 U758 ( .A(n4309), .B(n865), .C(n3846), .Y(n775) );
  AOI21X1 U760 ( .A(n809), .B(n4593), .C(n779), .Y(n777) );
  OAI21X1 U766 ( .A(n3215), .B(n2896), .C(n3087), .Y(n779) );
  XOR2X1 U771 ( .A(n3673), .B(n4085), .Y(SUM[124]) );
  AOI21X1 U772 ( .A(n4774), .B(n3086), .C(n788), .Y(n786) );
  OAI21X1 U774 ( .A(n3456), .B(n4793), .C(n3164), .Y(n788) );
  AOI21X1 U776 ( .A(n4719), .B(n4268), .C(n792), .Y(n790) );
  OAI21X1 U778 ( .A(n4308), .B(n865), .C(n3845), .Y(n792) );
  AOI21X1 U780 ( .A(n809), .B(n795), .C(n3748), .Y(n794) );
  XOR2X1 U787 ( .A(n3672), .B(n4084), .Y(SUM[123]) );
  AOI21X1 U788 ( .A(n4774), .B(n3085), .C(n801), .Y(n799) );
  OAI21X1 U790 ( .A(n3454), .B(n2874), .C(n3163), .Y(n801) );
  AOI21X1 U792 ( .A(n4753), .B(n4266), .C(n805), .Y(n803) );
  OAI21X1 U794 ( .A(n4688), .B(n865), .C(n4340), .Y(n805) );
  AOI21X1 U800 ( .A(n839), .B(n3254), .C(n813), .Y(n807) );
  OAI21X1 U802 ( .A(n4352), .B(n4502), .C(n3084), .Y(n813) );
  XOR2X1 U807 ( .A(n3671), .B(n4083), .Y(SUM[122]) );
  AOI21X1 U808 ( .A(n2865), .B(n2941), .C(n818), .Y(n816) );
  OAI21X1 U810 ( .A(n3453), .B(n2845), .C(n3162), .Y(n818) );
  AOI21X1 U812 ( .A(n4753), .B(n4264), .C(n822), .Y(n820) );
  OAI21X1 U814 ( .A(n4307), .B(n865), .C(n3844), .Y(n822) );
  AOI21X1 U816 ( .A(n839), .B(n827), .C(n828), .Y(n824) );
  XOR2X1 U823 ( .A(n3670), .B(n4082), .Y(SUM[121]) );
  AOI21X1 U824 ( .A(n4776), .B(n2940), .C(n831), .Y(n829) );
  OAI21X1 U826 ( .A(n3451), .B(n4793), .C(n3161), .Y(n831) );
  AOI21X1 U828 ( .A(n4753), .B(n4262), .C(n835), .Y(n833) );
  OAI21X1 U830 ( .A(n836), .B(n865), .C(n837), .Y(n835) );
  OAI21X1 U838 ( .A(n3480), .B(n4500), .C(n3083), .Y(n839) );
  XOR2X1 U843 ( .A(n3669), .B(n4081), .Y(SUM[120]) );
  AOI21X1 U844 ( .A(n4774), .B(n3082), .C(n848), .Y(n846) );
  OAI21X1 U846 ( .A(n3448), .B(n4793), .C(n3160), .Y(n848) );
  AOI21X1 U848 ( .A(n4753), .B(n4260), .C(n852), .Y(n850) );
  OAI21X1 U850 ( .A(n4603), .B(n865), .C(n4560), .Y(n852) );
  XOR2X1 U857 ( .A(n3668), .B(n4080), .Y(SUM[119]) );
  AOI21X1 U858 ( .A(n4659), .B(n3935), .C(n859), .Y(n857) );
  OAI21X1 U860 ( .A(n3447), .B(n2844), .C(n3843), .Y(n859) );
  AOI21X1 U862 ( .A(n4719), .B(n4636), .C(n863), .Y(n861) );
  OAI21X1 U868 ( .A(n3081), .B(n3536), .C(n3841), .Y(n863) );
  AOI21X1 U870 ( .A(n897), .B(n3080), .C(n871), .Y(n869) );
  OAI21X1 U872 ( .A(n4462), .B(n3518), .C(n3079), .Y(n871) );
  XOR2X1 U877 ( .A(n3667), .B(n4079), .Y(SUM[118]) );
  AOI21X1 U878 ( .A(n4774), .B(n3934), .C(n876), .Y(n874) );
  OAI21X1 U880 ( .A(n3445), .B(n4793), .C(n3839), .Y(n876) );
  AOI21X1 U882 ( .A(n4753), .B(n3078), .C(n880), .Y(n878) );
  OAI21X1 U884 ( .A(n4236), .B(n4390), .C(n4559), .Y(n880) );
  XOR2X1 U891 ( .A(n3666), .B(n4078), .Y(SUM[117]) );
  AOI21X1 U892 ( .A(n4774), .B(n2913), .C(n887), .Y(n885) );
  OAI21X1 U894 ( .A(n3443), .B(n4793), .C(n3837), .Y(n887) );
  AOI21X1 U896 ( .A(n4753), .B(n890), .C(n891), .Y(n889) );
  AOI21X1 U900 ( .A(n921), .B(n4538), .C(n897), .Y(n893) );
  OAI21X1 U904 ( .A(n3478), .B(n4249), .C(n3076), .Y(n897) );
  XOR2X1 U909 ( .A(n3665), .B(n4077), .Y(SUM[116]) );
  AOI21X1 U910 ( .A(n4776), .B(n2939), .C(n902), .Y(n900) );
  OAI21X1 U912 ( .A(n3442), .B(n4793), .C(n3835), .Y(n902) );
  AOI21X1 U914 ( .A(n4753), .B(n2938), .C(n906), .Y(n904) );
  OAI21X1 U916 ( .A(n4378), .B(n4582), .C(n3479), .Y(n906) );
  XOR2X1 U923 ( .A(n3664), .B(n4076), .Y(SUM[115]) );
  AOI21X1 U924 ( .A(n4774), .B(n2937), .C(n913), .Y(n911) );
  OAI21X1 U926 ( .A(n3440), .B(n4793), .C(n3833), .Y(n913) );
  AOI21X1 U928 ( .A(n4753), .B(n918), .C(n921), .Y(n915) );
  AOI21X1 U936 ( .A(n945), .B(n3318), .C(n925), .Y(n919) );
  OAI21X1 U938 ( .A(n4248), .B(n4461), .C(n3075), .Y(n925) );
  XOR2X1 U943 ( .A(n3663), .B(n4075), .Y(SUM[114]) );
  AOI21X1 U944 ( .A(n4774), .B(n2936), .C(n930), .Y(n928) );
  OAI21X1 U946 ( .A(n3438), .B(n4793), .C(n3831), .Y(n930) );
  AOI21X1 U948 ( .A(n4753), .B(n2935), .C(n934), .Y(n932) );
  OAI21X1 U950 ( .A(n4400), .B(n947), .C(n4558), .Y(n934) );
  XOR2X1 U957 ( .A(n3662), .B(n4074), .Y(SUM[113]) );
  AOI21X1 U958 ( .A(n4774), .B(n3074), .C(n941), .Y(n939) );
  OAI21X1 U960 ( .A(n3073), .B(n4793), .C(n3830), .Y(n941) );
  AOI21X1 U962 ( .A(n4718), .B(n4660), .C(n945), .Y(n943) );
  OAI21X1 U968 ( .A(n3214), .B(n3435), .C(n3072), .Y(n945) );
  XOR2X1 U973 ( .A(n3661), .B(n4073), .Y(SUM[112]) );
  AOI21X1 U974 ( .A(n4774), .B(n3071), .C(n954), .Y(n952) );
  OAI21X1 U976 ( .A(n3070), .B(n4793), .C(n3828), .Y(n954) );
  AOI21X1 U978 ( .A(n4753), .B(n959), .C(n3747), .Y(n956) );
  XOR2X1 U985 ( .A(n3660), .B(n4072), .Y(SUM[111]) );
  AOI21X1 U986 ( .A(n4774), .B(n3069), .C(n963), .Y(n961) );
  OAI21X1 U988 ( .A(n3326), .B(n4793), .C(n4722), .Y(n963) );
  AOI21X1 U994 ( .A(n1065), .B(n3729), .C(n971), .Y(n965) );
  OAI21X1 U996 ( .A(n3380), .B(n3535), .C(n3827), .Y(n971) );
  AOI21X1 U998 ( .A(n999), .B(n3068), .C(n975), .Y(n973) );
  OAI21X1 U1000 ( .A(n4350), .B(n3345), .C(n3067), .Y(n975) );
  XOR2X1 U1005 ( .A(n3659), .B(n4071), .Y(SUM[110]) );
  AOI21X1 U1006 ( .A(n4776), .B(n2934), .C(n980), .Y(n978) );
  OAI21X1 U1008 ( .A(n3066), .B(n2844), .C(n3825), .Y(n980) );
  AOI21X1 U1010 ( .A(n993), .B(n4184), .C(n984), .Y(n982) );
  XOR2X1 U1017 ( .A(n3658), .B(n4070), .Y(SUM[109]) );
  AOI21X1 U1018 ( .A(n4776), .B(n3065), .C(n989), .Y(n987) );
  OAI21X1 U1020 ( .A(n990), .B(n2844), .C(n991), .Y(n989) );
  OAI21X1 U1024 ( .A(n4306), .B(n1067), .C(n3824), .Y(n993) );
  AOI21X1 U1026 ( .A(n1021), .B(n4536), .C(n999), .Y(n995) );
  OAI21X1 U1030 ( .A(n4349), .B(n3978), .C(n3063), .Y(n999) );
  XOR2X1 U1035 ( .A(n3657), .B(n4069), .Y(SUM[108]) );
  AOI21X1 U1036 ( .A(n4776), .B(n3062), .C(n1004), .Y(n1002) );
  OAI21X1 U1038 ( .A(n3061), .B(n4793), .C(n3822), .Y(n1004) );
  AOI21X1 U1040 ( .A(n1017), .B(n1009), .C(n1010), .Y(n1006) );
  XOR2X1 U1047 ( .A(n3656), .B(n4068), .Y(SUM[107]) );
  AOI21X1 U1048 ( .A(n4775), .B(n3059), .C(n1013), .Y(n1011) );
  OAI21X1 U1054 ( .A(n4579), .B(n1067), .C(n4338), .Y(n1017) );
  AOI21X1 U1060 ( .A(n1047), .B(n4284), .C(n1025), .Y(n1019) );
  OAI21X1 U1062 ( .A(n4348), .B(n4496), .C(n3058), .Y(n1025) );
  XOR2X1 U1067 ( .A(n3655), .B(n4067), .Y(SUM[106]) );
  AOI21X1 U1068 ( .A(n4776), .B(n3057), .C(n1030), .Y(n1028) );
  OAI21X1 U1070 ( .A(n3056), .B(n4793), .C(n3820), .Y(n1030) );
  AOI21X1 U1072 ( .A(n1043), .B(n2181), .C(n1036), .Y(n1032) );
  XOR2X1 U1079 ( .A(n3654), .B(n4066), .Y(SUM[105]) );
  AOI21X1 U1080 ( .A(n4775), .B(n3055), .C(n1039), .Y(n1037) );
  OAI21X1 U1082 ( .A(n1040), .B(n4793), .C(n1041), .Y(n1039) );
  OAI21X1 U1086 ( .A(n1044), .B(n1067), .C(n1045), .Y(n1043) );
  OAI21X1 U1090 ( .A(n3213), .B(n4494), .C(n4203), .Y(n1047) );
  XOR2X1 U1095 ( .A(n3653), .B(n4065), .Y(SUM[104]) );
  AOI21X1 U1096 ( .A(n4774), .B(n3054), .C(n1052), .Y(n1050) );
  OAI21X1 U1098 ( .A(n4305), .B(n4793), .C(n3819), .Y(n1052) );
  AOI21X1 U1100 ( .A(n2893), .B(n3752), .C(n3746), .Y(n1054) );
  XOR2X1 U1107 ( .A(n3652), .B(n4064), .Y(SUM[103]) );
  AOI21X1 U1108 ( .A(n4776), .B(n3053), .C(n1061), .Y(n1059) );
  OAI21X1 U1110 ( .A(n2845), .B(n1064), .C(n1067), .Y(n1061) );
  OAI21X1 U1118 ( .A(n3595), .B(n3534), .C(n3159), .Y(n1065) );
  AOI21X1 U1120 ( .A(n1095), .B(n4282), .C(n1073), .Y(n1071) );
  OAI21X1 U1122 ( .A(n4346), .B(n3434), .C(n3050), .Y(n1073) );
  XOR2X1 U1127 ( .A(n3651), .B(n4063), .Y(SUM[102]) );
  AOI21X1 U1128 ( .A(n4775), .B(n2933), .C(n1078), .Y(n1076) );
  OAI21X1 U1130 ( .A(n4304), .B(n4793), .C(n3818), .Y(n1078) );
  AOI21X1 U1132 ( .A(n1091), .B(n4181), .C(n1082), .Y(n1080) );
  XOR2X1 U1139 ( .A(n3650), .B(n4062), .Y(SUM[101]) );
  AOI21X1 U1140 ( .A(n4775), .B(n3933), .C(n1087), .Y(n1085) );
  OAI21X1 U1142 ( .A(n1088), .B(n4793), .C(n1089), .Y(n1087) );
  OAI21X1 U1146 ( .A(n1092), .B(n3534), .C(n1093), .Y(n1091) );
  OAI21X1 U1150 ( .A(n3898), .B(n4493), .C(n3049), .Y(n1095) );
  XOR2X1 U1155 ( .A(n3649), .B(n4061), .Y(SUM[100]) );
  AOI21X1 U1156 ( .A(n4776), .B(n3048), .C(n1100), .Y(n1098) );
  OAI21X1 U1158 ( .A(n4303), .B(n4793), .C(n3817), .Y(n1100) );
  AOI21X1 U1160 ( .A(n1113), .B(n2187), .C(n4345), .Y(n1102) );
  XOR2X1 U1167 ( .A(n3648), .B(n4060), .Y(SUM[99]) );
  AOI21X1 U1168 ( .A(n4775), .B(n3047), .C(n1109), .Y(n1107) );
  OAI21X1 U1170 ( .A(n4723), .B(n4793), .C(n3534), .Y(n1109) );
  AOI21X1 U1180 ( .A(n1139), .B(n3559), .C(n1121), .Y(n1115) );
  OAI21X1 U1182 ( .A(n3466), .B(n4492), .C(n3045), .Y(n1121) );
  AOI21X1 U1188 ( .A(n4776), .B(n3044), .C(n1126), .Y(n1124) );
  OAI21X1 U1190 ( .A(n4302), .B(n4793), .C(n3816), .Y(n1126) );
  AOI21X1 U1192 ( .A(n2847), .B(n2189), .C(n1130), .Y(n1128) );
  XOR2X1 U1199 ( .A(n3647), .B(n4059), .Y(SUM[97]) );
  AOI21X1 U1200 ( .A(n4776), .B(n1134), .C(n1135), .Y(n1133) );
  OAI21X1 U1202 ( .A(n1136), .B(n2874), .C(n1137), .Y(n1135) );
  OAI21X1 U1210 ( .A(n4491), .B(n3220), .C(n3042), .Y(n1139) );
  XOR2X1 U1215 ( .A(n3646), .B(n4058), .Y(SUM[96]) );
  AOI21X1 U1216 ( .A(n4776), .B(n3041), .C(n1148), .Y(n1146) );
  OAI21X1 U1218 ( .A(n4601), .B(n4793), .C(n3220), .Y(n1148) );
  XOR2X1 U1225 ( .A(n3645), .B(n4057), .Y(SUM[95]) );
  AOI21X1 U1226 ( .A(n4776), .B(n4764), .C(n2875), .Y(n1153) );
  OAI21X1 U1232 ( .A(n2894), .B(n3505), .C(n3158), .Y(n1155) );
  AOI21X1 U1234 ( .A(n1249), .B(n3314), .C(n1163), .Y(n1161) );
  OAI21X1 U1236 ( .A(n3040), .B(n3533), .C(n3157), .Y(n1163) );
  AOI21X1 U1238 ( .A(n1189), .B(n3312), .C(n1167), .Y(n1165) );
  OAI21X1 U1240 ( .A(n4216), .B(n4246), .C(n3039), .Y(n1167) );
  XOR2X1 U1245 ( .A(n3644), .B(n4056), .Y(SUM[94]) );
  AOI21X1 U1246 ( .A(n4774), .B(n3038), .C(n1172), .Y(n1170) );
  OAI21X1 U1248 ( .A(n3204), .B(n4734), .C(n2955), .Y(n1172) );
  XOR2X1 U1255 ( .A(n3643), .B(n4055), .Y(SUM[93]) );
  AOI21X1 U1256 ( .A(n4659), .B(n1178), .C(n1179), .Y(n1177) );
  OAI21X1 U1262 ( .A(n4301), .B(n1251), .C(n3815), .Y(n1183) );
  AOI21X1 U1264 ( .A(n1209), .B(n3292), .C(n1189), .Y(n1185) );
  OAI21X1 U1268 ( .A(n2931), .B(n2914), .C(n4202), .Y(n1189) );
  XOR2X1 U1273 ( .A(n3642), .B(n4054), .Y(SUM[92]) );
  AOI21X1 U1274 ( .A(n4774), .B(n3037), .C(n1194), .Y(n1192) );
  OAI21X1 U1276 ( .A(n4234), .B(n4437), .C(n2931), .Y(n1194) );
  XOR2X1 U1283 ( .A(n3641), .B(n4053), .Y(SUM[91]) );
  AOI21X1 U1284 ( .A(n2865), .B(n1200), .C(n1201), .Y(n1199) );
  AOI21X1 U1288 ( .A(n1335), .B(n2930), .C(n1205), .Y(n1203) );
  OAI21X1 U1290 ( .A(n4772), .B(n1251), .C(n4337), .Y(n1205) );
  AOI21X1 U1296 ( .A(n1233), .B(n3036), .C(n1213), .Y(n1207) );
  OAI21X1 U1298 ( .A(n4245), .B(n4460), .C(n3035), .Y(n1213) );
  XOR2X1 U1303 ( .A(n3640), .B(n4052), .Y(SUM[90]) );
  AOI21X1 U1304 ( .A(n4774), .B(n3034), .C(n1218), .Y(n1216) );
  OAI21X1 U1306 ( .A(n3884), .B(n4729), .C(n3033), .Y(n1218) );
  XOR2X1 U1313 ( .A(n3639), .B(n4051), .Y(SUM[89]) );
  AOI21X1 U1314 ( .A(n4776), .B(n1224), .C(n1225), .Y(n1223) );
  AOI21X1 U1318 ( .A(n1335), .B(n2929), .C(n1229), .Y(n1227) );
  OAI21X1 U1320 ( .A(n1230), .B(n1251), .C(n1231), .Y(n1229) );
  OAI21X1 U1324 ( .A(n3476), .B(n4490), .C(n4201), .Y(n1233) );
  XOR2X1 U1329 ( .A(n3638), .B(n4050), .Y(SUM[88]) );
  AOI21X1 U1330 ( .A(n4775), .B(n3932), .C(n1238), .Y(n1236) );
  OAI21X1 U1332 ( .A(n3883), .B(n4407), .C(n4557), .Y(n1238) );
  XOR2X1 U1339 ( .A(n3637), .B(n4049), .Y(SUM[87]) );
  AOI21X1 U1340 ( .A(n4775), .B(n1244), .C(n1245), .Y(n1243) );
  AOI21X1 U1344 ( .A(n1335), .B(n4769), .C(n4669), .Y(n1247) );
  OAI21X1 U1350 ( .A(n3594), .B(n3532), .C(n3156), .Y(n1249) );
  AOI21X1 U1352 ( .A(n1277), .B(n3032), .C(n1257), .Y(n1255) );
  OAI21X1 U1354 ( .A(n4555), .B(n3031), .C(n4200), .Y(n1257) );
  XOR2X1 U1359 ( .A(n3636), .B(n4048), .Y(SUM[86]) );
  AOI21X1 U1360 ( .A(n4776), .B(n3931), .C(n1262), .Y(n1260) );
  OAI21X1 U1362 ( .A(n4233), .B(n4427), .C(n4556), .Y(n1262) );
  XOR2X1 U1369 ( .A(n3635), .B(n4047), .Y(SUM[85]) );
  AOI21X1 U1370 ( .A(n4775), .B(n1268), .C(n1269), .Y(n1267) );
  AOI21X1 U1374 ( .A(n1335), .B(n4281), .C(n1273), .Y(n1271) );
  OAI21X1 U1376 ( .A(n1274), .B(n3532), .C(n1275), .Y(n1273) );
  OAI21X1 U1380 ( .A(n3030), .B(n4489), .C(n4199), .Y(n1277) );
  XOR2X1 U1385 ( .A(n3634), .B(n4046), .Y(SUM[84]) );
  AOI21X1 U1386 ( .A(n4775), .B(n3930), .C(n1282), .Y(n1280) );
  OAI21X1 U1388 ( .A(n3882), .B(n4411), .C(n3030), .Y(n1282) );
  XOR2X1 U1395 ( .A(n3633), .B(n4045), .Y(SUM[83]) );
  AOI21X1 U1396 ( .A(n4776), .B(n1290), .C(n1289), .Y(n1287) );
  AOI21X1 U1400 ( .A(n1335), .B(n1292), .C(n1293), .Y(n1291) );
  AOI21X1 U1408 ( .A(n1319), .B(n3028), .C(n1301), .Y(n1295) );
  OAI21X1 U1410 ( .A(n2928), .B(n3400), .C(n4198), .Y(n1301) );
  XOR2X1 U1415 ( .A(n3632), .B(n4044), .Y(SUM[82]) );
  AOI21X1 U1416 ( .A(n4776), .B(n3929), .C(n1306), .Y(n1304) );
  OAI21X1 U1418 ( .A(n3881), .B(n4432), .C(n2928), .Y(n1306) );
  XOR2X1 U1425 ( .A(n3631), .B(n4043), .Y(SUM[81]) );
  AOI21X1 U1426 ( .A(n4775), .B(n1312), .C(n1313), .Y(n1311) );
  AOI21X1 U1430 ( .A(n1335), .B(n3290), .C(n1319), .Y(n1315) );
  OAI21X1 U1434 ( .A(n3474), .B(n4487), .C(n4197), .Y(n1319) );
  XOR2X1 U1439 ( .A(n3630), .B(n4042), .Y(SUM[80]) );
  AOI21X1 U1440 ( .A(n4659), .B(n3928), .C(n1324), .Y(n1322) );
  OAI21X1 U1442 ( .A(n4430), .B(n4786), .C(n3475), .Y(n1324) );
  XOR2X1 U1449 ( .A(n3629), .B(n4041), .Y(SUM[79]) );
  AOI21X1 U1450 ( .A(n4774), .B(n2848), .C(n1335), .Y(n1329) );
  AOI21X1 U1458 ( .A(n2881), .B(n2902), .C(n1339), .Y(n1333) );
  OAI21X1 U1460 ( .A(n4716), .B(n3504), .C(n3813), .Y(n1339) );
  AOI21X1 U1462 ( .A(n1361), .B(n3245), .C(n1343), .Y(n1341) );
  OAI21X1 U1464 ( .A(n4244), .B(n3343), .C(n4196), .Y(n1343) );
  XOR2X1 U1469 ( .A(n3628), .B(n4040), .Y(SUM[78]) );
  AOI21X1 U1470 ( .A(n4775), .B(n3927), .C(n1348), .Y(n1346) );
  OAI21X1 U1472 ( .A(n4664), .B(n3531), .C(n3027), .Y(n1348) );
  XOR2X1 U1479 ( .A(n3627), .B(n4039), .Y(SUM[77]) );
  AOI21X1 U1480 ( .A(n4775), .B(n1354), .C(n1355), .Y(n1353) );
  AOI21X1 U1484 ( .A(n1373), .B(n3266), .C(n1361), .Y(n1357) );
  OAI21X1 U1488 ( .A(n2871), .B(n3516), .C(n3026), .Y(n1361) );
  XOR2X1 U1493 ( .A(n3626), .B(n4038), .Y(SUM[76]) );
  AOI21X1 U1494 ( .A(n4775), .B(n3926), .C(n1366), .Y(n1364) );
  OAI21X1 U1496 ( .A(n4434), .B(n1375), .C(n4554), .Y(n1366) );
  XOR2X1 U1503 ( .A(n3625), .B(n4037), .Y(SUM[75]) );
  AOI21X1 U1504 ( .A(n4775), .B(n4328), .C(n1373), .Y(n1371) );
  OAI21X1 U1510 ( .A(n3325), .B(n4641), .C(n4289), .Y(n1373) );
  AOI21X1 U1514 ( .A(n1401), .B(n4280), .C(n1383), .Y(n1381) );
  OAI21X1 U1516 ( .A(n2922), .B(n4459), .C(n3024), .Y(n1383) );
  XOR2X1 U1521 ( .A(n3624), .B(n4036), .Y(SUM[74]) );
  AOI21X1 U1522 ( .A(n2865), .B(n3925), .C(n1388), .Y(n1386) );
  OAI21X1 U1524 ( .A(n4766), .B(n3530), .C(n4553), .Y(n1388) );
  XOR2X1 U1531 ( .A(n3623), .B(n4035), .Y(SUM[73]) );
  AOI21X1 U1532 ( .A(n4774), .B(n1394), .C(n1395), .Y(n1393) );
  AOI21X1 U1536 ( .A(n4642), .B(n4534), .C(n2892), .Y(n1397) );
  OAI21X1 U1540 ( .A(n3908), .B(n3219), .C(n3022), .Y(n1401) );
  XOR2X1 U1545 ( .A(n3622), .B(n4034), .Y(SUM[72]) );
  AOI21X1 U1546 ( .A(n4775), .B(n3924), .C(n1406), .Y(n1404) );
  OAI21X1 U1548 ( .A(n4756), .B(n4641), .C(n3219), .Y(n1406) );
  XOR2X1 U1555 ( .A(n3621), .B(n4033), .Y(SUM[71]) );
  AOI21X1 U1556 ( .A(n4776), .B(n2884), .C(n4642), .Y(n1411) );
  AOI21X1 U1568 ( .A(n4665), .B(n1443), .C(n1425), .Y(n1423) );
  OAI21X1 U1570 ( .A(n4457), .B(n3508), .C(n4195), .Y(n1425) );
  XOR2X1 U1575 ( .A(n3620), .B(n4032), .Y(SUM[70]) );
  AOI21X1 U1576 ( .A(n4776), .B(n3923), .C(n1430), .Y(n1428) );
  OAI21X1 U1578 ( .A(n4232), .B(n4441), .C(n3507), .Y(n1430) );
  XOR2X1 U1585 ( .A(n3619), .B(n4031), .Y(SUM[69]) );
  AOI21X1 U1586 ( .A(n4775), .B(n1436), .C(n1437), .Y(n1435) );
  AOI21X1 U1590 ( .A(n1459), .B(n3300), .C(n1443), .Y(n1439) );
  OAI21X1 U1594 ( .A(n2916), .B(n4485), .C(n4194), .Y(n1443) );
  XOR2X1 U1599 ( .A(n3618), .B(n4030), .Y(SUM[68]) );
  AOI21X1 U1600 ( .A(n4774), .B(n2927), .C(n1448), .Y(n1446) );
  OAI21X1 U1602 ( .A(n4445), .B(n4757), .C(n2916), .Y(n1448) );
  XOR2X1 U1609 ( .A(n3617), .B(n4029), .Y(SUM[67]) );
  AOI21X1 U1610 ( .A(n4774), .B(n4714), .C(n1459), .Y(n1453) );
  AOI21X1 U1618 ( .A(n1475), .B(n3250), .C(n1463), .Y(n1457) );
  OAI21X1 U1620 ( .A(n2921), .B(n4455), .C(n3020), .Y(n1463) );
  XOR2X1 U1625 ( .A(n3616), .B(n4028), .Y(SUM[66]) );
  AOI21X1 U1626 ( .A(n4775), .B(n3922), .C(n1468), .Y(n1466) );
  OAI21X1 U1628 ( .A(n4765), .B(n1477), .C(n2921), .Y(n1468) );
  XOR2X1 U1635 ( .A(n3615), .B(n4027), .Y(SUM[65]) );
  AOI21X1 U1636 ( .A(n4775), .B(n4707), .C(n2880), .Y(n1473) );
  OAI21X1 U1642 ( .A(n3472), .B(n3230), .C(n3019), .Y(n1475) );
  AOI21X1 U1648 ( .A(n4775), .B(n1485), .C(n1484), .Y(n1482) );
  XNOR2X1 U1655 ( .A(n1501), .B(n4014), .Y(SUM[63]) );
  AOI21X1 U1657 ( .A(n2860), .B(n3921), .C(n1490), .Y(n1488) );
  OAI21X1 U1659 ( .A(n3573), .B(n3527), .C(n3154), .Y(n1490) );
  AOI21X1 U1661 ( .A(n1594), .B(n4693), .C(n1494), .Y(n1492) );
  OAI21X1 U1663 ( .A(n3428), .B(n3529), .C(n3811), .Y(n1494) );
  AOI21X1 U1665 ( .A(n1522), .B(n3243), .C(n1498), .Y(n1496) );
  OAI21X1 U1667 ( .A(n4243), .B(n4454), .C(n3018), .Y(n1498) );
  XNOR2X1 U1672 ( .A(n1514), .B(n4013), .Y(SUM[62]) );
  OAI21X1 U1673 ( .A(n3975), .B(n2911), .C(n3809), .Y(n1501) );
  AOI21X1 U1675 ( .A(n1682), .B(n2901), .C(n1505), .Y(n1503) );
  OAI21X1 U1677 ( .A(n4300), .B(n1596), .C(n3807), .Y(n1505) );
  AOI21X1 U1679 ( .A(n1548), .B(n4254), .C(n1509), .Y(n1507) );
  OAI21X1 U1681 ( .A(n4730), .B(n1524), .C(n4552), .Y(n1509) );
  XNOR2X1 U1688 ( .A(n1529), .B(n4012), .Y(SUM[61]) );
  OAI21X1 U1689 ( .A(n3974), .B(n3740), .C(n3806), .Y(n1514) );
  AOI21X1 U1691 ( .A(n1682), .B(n3016), .C(n1518), .Y(n1516) );
  OAI21X1 U1693 ( .A(n4299), .B(n1596), .C(n3804), .Y(n1518) );
  AOI21X1 U1695 ( .A(n1548), .B(n4710), .C(n1522), .Y(n1520) );
  OAI21X1 U1701 ( .A(n3212), .B(n4483), .C(n3014), .Y(n1522) );
  XNOR2X1 U1706 ( .A(n1540), .B(n4011), .Y(SUM[60]) );
  OAI21X1 U1707 ( .A(n3973), .B(n4794), .C(n3803), .Y(n1529) );
  AOI21X1 U1709 ( .A(n1682), .B(n3013), .C(n1533), .Y(n1531) );
  OAI21X1 U1711 ( .A(n4298), .B(n1596), .C(n3801), .Y(n1533) );
  AOI21X1 U1713 ( .A(n1548), .B(n2227), .C(n1539), .Y(n1535) );
  XNOR2X1 U1720 ( .A(n1555), .B(n4010), .Y(SUM[59]) );
  OAI21X1 U1721 ( .A(n3972), .B(n4794), .C(n3800), .Y(n1540) );
  AOI21X1 U1723 ( .A(n1682), .B(n3012), .C(n1544), .Y(n1542) );
  OAI21X1 U1725 ( .A(n4742), .B(n1596), .C(n4336), .Y(n1544) );
  AOI21X1 U1731 ( .A(n1574), .B(n3241), .C(n1552), .Y(n1546) );
  OAI21X1 U1733 ( .A(n3211), .B(n4482), .C(n3011), .Y(n1552) );
  XNOR2X1 U1738 ( .A(n1566), .B(n4009), .Y(SUM[58]) );
  OAI21X1 U1739 ( .A(n3971), .B(n4794), .C(n3798), .Y(n1555) );
  AOI21X1 U1741 ( .A(n1682), .B(n3010), .C(n1559), .Y(n1557) );
  OAI21X1 U1743 ( .A(n4297), .B(n1596), .C(n3796), .Y(n1559) );
  AOI21X1 U1745 ( .A(n1574), .B(n2229), .C(n3745), .Y(n1561) );
  XNOR2X1 U1752 ( .A(n1581), .B(n4008), .Y(SUM[57]) );
  OAI21X1 U1753 ( .A(n3970), .B(n4794), .C(n3795), .Y(n1566) );
  AOI21X1 U1755 ( .A(n1682), .B(n3009), .C(n1570), .Y(n1568) );
  OAI21X1 U1757 ( .A(n1571), .B(n1596), .C(n1572), .Y(n1570) );
  OAI21X1 U1765 ( .A(n2920), .B(n4452), .C(n3008), .Y(n1574) );
  OAI21X1 U1771 ( .A(n3969), .B(n2911), .C(n3793), .Y(n1581) );
  AOI21X1 U1773 ( .A(n1682), .B(n3007), .C(n1585), .Y(n1583) );
  OAI21X1 U1775 ( .A(n4711), .B(n1596), .C(n2920), .Y(n1585) );
  XNOR2X1 U1782 ( .A(n1605), .B(n4006), .Y(SUM[55]) );
  OAI21X1 U1783 ( .A(n3968), .B(n4794), .C(n3791), .Y(n1590) );
  AOI21X1 U1785 ( .A(n1682), .B(n4739), .C(n4731), .Y(n1592) );
  OAI21X1 U1791 ( .A(n3424), .B(n3528), .C(n3789), .Y(n1594) );
  AOI21X1 U1793 ( .A(n1624), .B(n3006), .C(n1602), .Y(n1600) );
  OAI21X1 U1795 ( .A(n2919), .B(n4451), .C(n3004), .Y(n1602) );
  XNOR2X1 U1800 ( .A(n1614), .B(n4005), .Y(SUM[54]) );
  OAI21X1 U1801 ( .A(n3967), .B(n4794), .C(n3787), .Y(n1605) );
  AOI21X1 U1803 ( .A(n1682), .B(n4278), .C(n1609), .Y(n1607) );
  OAI21X1 U1805 ( .A(n4231), .B(n4721), .C(n2919), .Y(n1609) );
  XNOR2X1 U1812 ( .A(n1627), .B(n4004), .Y(SUM[53]) );
  OAI21X1 U1813 ( .A(n3966), .B(n4794), .C(n3785), .Y(n1614) );
  AOI21X1 U1815 ( .A(n1682), .B(n1617), .C(n1618), .Y(n1616) );
  AOI21X1 U1819 ( .A(n4580), .B(n4532), .C(n1624), .Y(n1620) );
  OAI21X1 U1823 ( .A(n4360), .B(n3229), .C(n3003), .Y(n1624) );
  OAI21X1 U1829 ( .A(n3965), .B(n4794), .C(n3783), .Y(n1627) );
  AOI21X1 U1831 ( .A(n1682), .B(n2925), .C(n1631), .Y(n1629) );
  OAI21X1 U1833 ( .A(n4703), .B(n4581), .C(n4361), .Y(n1631) );
  XNOR2X1 U1840 ( .A(n1651), .B(n4003), .Y(SUM[51]) );
  OAI21X1 U1841 ( .A(n3964), .B(n4794), .C(n3781), .Y(n1636) );
  AOI21X1 U1843 ( .A(n1682), .B(n2861), .C(n4580), .Y(n1638) );
  AOI21X1 U1851 ( .A(n1664), .B(n4277), .C(n1648), .Y(n1642) );
  OAI21X1 U1853 ( .A(n3468), .B(n4450), .C(n3002), .Y(n1648) );
  OAI21X1 U1859 ( .A(n3963), .B(n3740), .C(n3779), .Y(n1651) );
  AOI21X1 U1861 ( .A(n1682), .B(n4276), .C(n1655), .Y(n1653) );
  OAI21X1 U1863 ( .A(n4668), .B(n1666), .C(n4551), .Y(n1655) );
  XNOR2X1 U1870 ( .A(n1671), .B(n4002), .Y(SUM[49]) );
  OAI21X1 U1871 ( .A(n3962), .B(n2911), .C(n3777), .Y(n1660) );
  AOI21X1 U1873 ( .A(n1682), .B(n4592), .C(n1664), .Y(n1662) );
  OAI21X1 U1879 ( .A(n3870), .B(n3897), .C(n3001), .Y(n1664) );
  XNOR2X1 U1884 ( .A(n1678), .B(n4001), .Y(SUM[48]) );
  OAI21X1 U1885 ( .A(n3961), .B(n4794), .C(n3775), .Y(n1671) );
  AOI21X1 U1887 ( .A(n1682), .B(n1676), .C(n3744), .Y(n1673) );
  XNOR2X1 U1894 ( .A(n1693), .B(n4000), .Y(SUM[47]) );
  OAI21X1 U1895 ( .A(n4640), .B(n4794), .C(n4709), .Y(n1678) );
  AOI21X1 U1901 ( .A(n1764), .B(n2912), .C(n1686), .Y(n1680) );
  OAI21X1 U1903 ( .A(n3370), .B(n3526), .C(n3153), .Y(n1686) );
  AOI21X1 U1905 ( .A(n1710), .B(n3264), .C(n1690), .Y(n1688) );
  OAI21X1 U1907 ( .A(n4479), .B(n4356), .C(n3000), .Y(n1690) );
  XNOR2X1 U1912 ( .A(n1700), .B(n3999), .Y(SUM[46]) );
  OAI21X1 U1913 ( .A(n3960), .B(n4794), .C(n3773), .Y(n1693) );
  AOI21X1 U1915 ( .A(n1704), .B(n4149), .C(n1697), .Y(n1695) );
  XNOR2X1 U1922 ( .A(n1713), .B(n3998), .Y(SUM[45]) );
  OAI21X1 U1923 ( .A(n1701), .B(n4794), .C(n1702), .Y(n1700) );
  OAI21X1 U1927 ( .A(n4296), .B(n4643), .C(n3772), .Y(n1704) );
  AOI21X1 U1929 ( .A(n1728), .B(n3248), .C(n1710), .Y(n1706) );
  OAI21X1 U1933 ( .A(n3406), .B(n4325), .C(n2998), .Y(n1710) );
  OAI21X1 U1939 ( .A(n3959), .B(n3740), .C(n3771), .Y(n1713) );
  AOI21X1 U1941 ( .A(n1724), .B(n4170), .C(n1717), .Y(n1715) );
  XNOR2X1 U1948 ( .A(n1735), .B(n3997), .Y(SUM[43]) );
  OAI21X1 U1949 ( .A(n1721), .B(n2911), .C(n1722), .Y(n1720) );
  OAI21X1 U1953 ( .A(n4699), .B(n4643), .C(n4335), .Y(n1724) );
  AOI21X1 U1959 ( .A(n1750), .B(n3557), .C(n1732), .Y(n1726) );
  OAI21X1 U1961 ( .A(n3499), .B(n4478), .C(n2995), .Y(n1732) );
  XNOR2X1 U1966 ( .A(n1742), .B(n3996), .Y(SUM[42]) );
  OAI21X1 U1967 ( .A(n3958), .B(n4794), .C(n3770), .Y(n1735) );
  AOI21X1 U1969 ( .A(n1746), .B(n1740), .C(n1741), .Y(n1737) );
  XNOR2X1 U1976 ( .A(n1753), .B(n3995), .Y(SUM[41]) );
  OAI21X1 U1977 ( .A(n1743), .B(n4794), .C(n1744), .Y(n1742) );
  OAI21X1 U1981 ( .A(n1747), .B(n4643), .C(n1748), .Y(n1746) );
  OAI21X1 U1985 ( .A(n2856), .B(n3223), .C(n2994), .Y(n1750) );
  XNOR2X1 U1990 ( .A(n1760), .B(n3994), .Y(SUM[40]) );
  OAI21X1 U1991 ( .A(n3957), .B(n4794), .C(n3769), .Y(n1753) );
  AOI21X1 U1993 ( .A(n2898), .B(n1758), .C(n3750), .Y(n1755) );
  XNOR2X1 U2000 ( .A(n1775), .B(n3993), .Y(SUM[39]) );
  OAI21X1 U2001 ( .A(n1765), .B(n4794), .C(n4643), .Y(n1760) );
  OAI21X1 U2009 ( .A(n2993), .B(n3502), .C(n3152), .Y(n1764) );
  AOI21X1 U2011 ( .A(n1790), .B(n2859), .C(n1772), .Y(n1770) );
  OAI21X1 U2013 ( .A(n3420), .B(n4355), .C(n2992), .Y(n1772) );
  XNOR2X1 U2018 ( .A(n1782), .B(n3992), .Y(SUM[38]) );
  OAI21X1 U2019 ( .A(n3956), .B(n2911), .C(n3768), .Y(n1775) );
  AOI21X1 U2021 ( .A(n1786), .B(n2891), .C(n1779), .Y(n1777) );
  XNOR2X1 U2028 ( .A(n1793), .B(n3991), .Y(SUM[37]) );
  OAI21X1 U2029 ( .A(n1783), .B(n3740), .C(n1784), .Y(n1782) );
  OAI21X1 U2033 ( .A(n1787), .B(n4767), .C(n1788), .Y(n1786) );
  OAI21X1 U2037 ( .A(n4344), .B(n4476), .C(n4193), .Y(n1790) );
  XNOR2X1 U2042 ( .A(n1800), .B(n3990), .Y(SUM[36]) );
  OAI21X1 U2043 ( .A(n3955), .B(n4794), .C(n3767), .Y(n1793) );
  AOI21X1 U2045 ( .A(n1804), .B(n2251), .C(n1797), .Y(n1795) );
  XNOR2X1 U2052 ( .A(n1815), .B(n3989), .Y(SUM[35]) );
  OAI21X1 U2053 ( .A(n3335), .B(n4794), .C(n4767), .Y(n1800) );
  AOI21X1 U2063 ( .A(n1826), .B(n3568), .C(n1812), .Y(n1806) );
  OAI21X1 U2065 ( .A(n3592), .B(n3556), .C(n2989), .Y(n1812) );
  XNOR2X1 U2070 ( .A(n1822), .B(n3988), .Y(SUM[34]) );
  OAI21X1 U2071 ( .A(n3954), .B(n4794), .C(n3766), .Y(n1815) );
  AOI21X1 U2073 ( .A(n2897), .B(n2253), .C(n1819), .Y(n1817) );
  XNOR2X1 U2080 ( .A(n1833), .B(n3987), .Y(SUM[33]) );
  OAI21X1 U2081 ( .A(n1823), .B(n4794), .C(n1824), .Y(n1822) );
  OAI21X1 U2089 ( .A(n3880), .B(n3514), .C(n3288), .Y(n1826) );
  OAI21X1 U2095 ( .A(n4358), .B(n2911), .C(n3513), .Y(n1833) );
  XOR2X1 U2100 ( .A(n3980), .B(n4026), .Y(SUM[31]) );
  AOI21X1 U2104 ( .A(n2867), .B(n1925), .C(n1841), .Y(n1839) );
  OAI21X1 U2106 ( .A(n3416), .B(n4333), .C(n3150), .Y(n1841) );
  AOI21X1 U2108 ( .A(n1865), .B(n3240), .C(n1845), .Y(n1843) );
  OAI21X1 U2110 ( .A(n2985), .B(n3888), .C(n2987), .Y(n1845) );
  XOR2X1 U2115 ( .A(n3614), .B(n4025), .Y(SUM[30]) );
  AOI21X1 U2116 ( .A(n2837), .B(n2986), .C(n1850), .Y(n1848) );
  OAI21X1 U2118 ( .A(n4295), .B(n1927), .C(n3765), .Y(n1850) );
  AOI21X1 U2120 ( .A(n1887), .B(n3261), .C(n1854), .Y(n1852) );
  OAI21X1 U2122 ( .A(n4424), .B(n1867), .C(n2985), .Y(n1854) );
  XOR2X1 U2129 ( .A(n3613), .B(n4024), .Y(SUM[29]) );
  AOI21X1 U2130 ( .A(n2836), .B(n2984), .C(n1861), .Y(n1859) );
  OAI21X1 U2132 ( .A(n4294), .B(n1927), .C(n3764), .Y(n1861) );
  AOI21X1 U2134 ( .A(n1887), .B(n4701), .C(n1865), .Y(n1863) );
  OAI21X1 U2140 ( .A(n3210), .B(n4475), .C(n2981), .Y(n1865) );
  XOR2X1 U2145 ( .A(n3612), .B(n4023), .Y(SUM[28]) );
  AOI21X1 U2146 ( .A(n4727), .B(n2980), .C(n1874), .Y(n1872) );
  OAI21X1 U2148 ( .A(n4293), .B(n1927), .C(n3763), .Y(n1874) );
  AOI21X1 U2150 ( .A(n1887), .B(n4148), .C(n1880), .Y(n1876) );
  AOI21X1 U2158 ( .A(n4727), .B(n2979), .C(n1883), .Y(n1881) );
  OAI21X1 U2160 ( .A(n4752), .B(n1927), .C(n4333), .Y(n1883) );
  AOI21X1 U2166 ( .A(n1909), .B(n4275), .C(n1891), .Y(n1885) );
  OAI21X1 U2168 ( .A(n4322), .B(n3404), .C(n2977), .Y(n1891) );
  AOI21X1 U2174 ( .A(n2837), .B(n2976), .C(n1896), .Y(n1894) );
  OAI21X1 U2176 ( .A(n4292), .B(n1927), .C(n3762), .Y(n1896) );
  AOI21X1 U2178 ( .A(n1909), .B(n4168), .C(n1900), .Y(n1898) );
  XOR2X1 U2185 ( .A(n3611), .B(n2924), .Y(SUM[25]) );
  AOI21X1 U2186 ( .A(n2836), .B(n2974), .C(n1905), .Y(n1903) );
  OAI21X1 U2188 ( .A(n1906), .B(n1927), .C(n1907), .Y(n1905) );
  OAI21X1 U2196 ( .A(n3209), .B(n3227), .C(n2973), .Y(n1909) );
  XOR2X1 U2201 ( .A(n3610), .B(n4022), .Y(SUM[24]) );
  AOI21X1 U2202 ( .A(n4727), .B(n2972), .C(n1918), .Y(n1916) );
  OAI21X1 U2204 ( .A(n4661), .B(n1927), .C(n3209), .Y(n1918) );
  XOR2X1 U2211 ( .A(n3609), .B(n4021), .Y(SUM[23]) );
  AOI21X1 U2212 ( .A(n2836), .B(n4635), .C(n4667), .Y(n1923) );
  OAI21X1 U2218 ( .A(n3498), .B(n3525), .C(n3149), .Y(n1925) );
  AOI21X1 U2220 ( .A(n3566), .B(n1951), .C(n1933), .Y(n1931) );
  OAI21X1 U2222 ( .A(n4359), .B(n4474), .C(n4192), .Y(n1933) );
  AOI21X1 U2228 ( .A(n4727), .B(n3920), .C(n1938), .Y(n1936) );
  OAI21X1 U2230 ( .A(n4230), .B(n4733), .C(n2970), .Y(n1938) );
  XOR2X1 U2237 ( .A(n3608), .B(n4020), .Y(SUM[21]) );
  AOI21X1 U2238 ( .A(n4727), .B(n4145), .C(n1945), .Y(n1943) );
  AOI21X1 U2242 ( .A(n1967), .B(n3238), .C(n1951), .Y(n1947) );
  OAI21X1 U2246 ( .A(n2915), .B(n3221), .C(n2969), .Y(n1951) );
  XOR2X1 U2251 ( .A(n3607), .B(n4019), .Y(SUM[20]) );
  AOI21X1 U2252 ( .A(n2837), .B(n3919), .C(n1956), .Y(n1954) );
  OAI21X1 U2254 ( .A(n4751), .B(n4726), .C(n4550), .Y(n1956) );
  XOR2X1 U2261 ( .A(n1974), .B(n4018), .Y(SUM[19]) );
  AOI21X1 U2262 ( .A(n2837), .B(n1966), .C(n1967), .Y(n1961) );
  AOI21X1 U2270 ( .A(n1983), .B(n4210), .C(n1971), .Y(n1965) );
  OAI21X1 U2272 ( .A(n2966), .B(n4472), .C(n2967), .Y(n1971) );
  OAI21X1 U2280 ( .A(n4780), .B(n1985), .C(n2966), .Y(n1976) );
  XOR2X1 U2287 ( .A(n3606), .B(n4017), .Y(SUM[17]) );
  OAI21X1 U2294 ( .A(n3408), .B(n3226), .C(n2965), .Y(n1983) );
  AOI21X1 U2300 ( .A(n2836), .B(n1993), .C(n3743), .Y(n1990) );
  XNOR2X1 U2307 ( .A(n2005), .B(n3986), .Y(SUM[15]) );
  AOI21X1 U2309 ( .A(n2065), .B(n3918), .C(n1998), .Y(n1996) );
  OAI21X1 U2311 ( .A(n3590), .B(n3501), .C(n3148), .Y(n1998) );
  AOI21X1 U2313 ( .A(n2018), .B(n3236), .C(n2002), .Y(n2000) );
  OAI21X1 U2315 ( .A(n2964), .B(n3512), .C(n4191), .Y(n2002) );
  XNOR2X1 U2320 ( .A(n2014), .B(n3985), .Y(SUM[14]) );
  OAI21X1 U2321 ( .A(n3953), .B(n2064), .C(n3761), .Y(n2005) );
  AOI21X1 U2323 ( .A(n2036), .B(n4258), .C(n2009), .Y(n2007) );
  OAI21X1 U2325 ( .A(n4404), .B(n2020), .C(n3511), .Y(n2009) );
  XNOR2X1 U2332 ( .A(n2025), .B(n3984), .Y(SUM[13]) );
  OAI21X1 U2333 ( .A(n3952), .B(n2064), .C(n3759), .Y(n2014) );
  AOI21X1 U2335 ( .A(n2036), .B(n4763), .C(n2018), .Y(n2016) );
  OAI21X1 U2341 ( .A(n3208), .B(n3979), .C(n4190), .Y(n2018) );
  XNOR2X1 U2346 ( .A(n2032), .B(n3983), .Y(SUM[12]) );
  OAI21X1 U2347 ( .A(n3951), .B(n2064), .C(n3757), .Y(n2025) );
  AOI21X1 U2349 ( .A(n2036), .B(n2275), .C(n3742), .Y(n2027) );
  XNOR2X1 U2356 ( .A(n2043), .B(n3982), .Y(SUM[11]) );
  OAI21X1 U2357 ( .A(n3885), .B(n2064), .C(n4680), .Y(n2032) );
  AOI21X1 U2363 ( .A(n2054), .B(n2862), .C(n2040), .Y(n2034) );
  OAI21X1 U2365 ( .A(n3588), .B(n3510), .C(n2963), .Y(n2040) );
  OAI21X1 U2371 ( .A(n3950), .B(n2064), .C(n3755), .Y(n2043) );
  AOI21X1 U2373 ( .A(n2054), .B(n2048), .C(n4678), .Y(n2045) );
  XNOR2X1 U2380 ( .A(n2061), .B(n3981), .Y(SUM[9]) );
  OAI21X1 U2381 ( .A(n2051), .B(n2064), .C(n2052), .Y(n2050) );
  OAI21X1 U2389 ( .A(n3496), .B(n3222), .C(n2962), .Y(n2054) );
  OAI21X1 U2395 ( .A(n4357), .B(n2064), .C(n3497), .Y(n2061) );
  OAI21X1 U2402 ( .A(n3207), .B(n3500), .C(n3147), .Y(n2065) );
  AOI21X1 U2404 ( .A(n3316), .B(n2081), .C(n2069), .Y(n2067) );
  OAI21X1 U2406 ( .A(n2959), .B(n3224), .C(n2960), .Y(n2069) );
  XOR2X1 U2411 ( .A(n3605), .B(n4016), .Y(SUM[6]) );
  OAI21X1 U2414 ( .A(n2075), .B(n2083), .C(n2959), .Y(n2074) );
  AOI21X1 U2422 ( .A(n2093), .B(n4326), .C(n2081), .Y(n2079) );
  OAI21X1 U2428 ( .A(n3206), .B(n3225), .C(n2958), .Y(n2081) );
  AOI21X1 U2434 ( .A(n2093), .B(n2091), .C(n3892), .Y(n2088) );
  AOI21X1 U2443 ( .A(n2103), .B(n3203), .C(n2096), .Y(n2094) );
  OAI21X1 U2445 ( .A(n3494), .B(n3603), .C(n2957), .Y(n2096) );
  XOR2X1 U2450 ( .A(n2102), .B(n3732), .Y(SUM[2]) );
  OAI21X1 U2451 ( .A(n4639), .B(n2102), .C(n3495), .Y(n2099) );
  OAI21X1 U2458 ( .A(n3205), .B(n2854), .C(n2956), .Y(n2103) );
  INVX4 U2471 ( .A(n2851), .Y(n2064) );
  OAI21X1 U2472 ( .A(n4662), .B(n1975), .C(n2835), .Y(n2834) );
  INVX2 U2473 ( .A(n2834), .Y(n1974) );
  INVX8 U2474 ( .A(n1976), .Y(n2835) );
  INVX2 U2475 ( .A(n4662), .Y(n2836) );
  INVX2 U2476 ( .A(n4662), .Y(n2837) );
  INVX2 U2477 ( .A(n4662), .Y(n4727) );
  XNOR2X1 U2478 ( .A(n2838), .B(n133), .Y(SUM[64]) );
  INVX1 U2479 ( .A(n2865), .Y(n2838) );
  OAI21X1 U2480 ( .A(n3123), .B(n3540), .C(n3168), .Y(n2839) );
  AND2X2 U2481 ( .A(n4179), .B(n4180), .Y(n2840) );
  INVX1 U2482 ( .A(n1064), .Y(n2841) );
  INVX1 U2483 ( .A(n1064), .Y(n2842) );
  OAI21X1 U2484 ( .A(n4217), .B(n3503), .C(n3155), .Y(n2843) );
  INVX1 U2485 ( .A(n4787), .Y(n2844) );
  INVX1 U2486 ( .A(n4787), .Y(n2845) );
  AND2X2 U2487 ( .A(n918), .B(n868), .Y(n2846) );
  INVX4 U2488 ( .A(n2846), .Y(n862) );
  INVX1 U2489 ( .A(n1137), .Y(n2847) );
  AND2X2 U2490 ( .A(n4141), .B(n2884), .Y(n2848) );
  AND2X2 U2491 ( .A(n1160), .B(n1332), .Y(n2849) );
  AND2X2 U2492 ( .A(n1160), .B(n1332), .Y(n2850) );
  OAI21X1 U2493 ( .A(n3207), .B(n3500), .C(n3147), .Y(n2851) );
  AND2X2 U2494 ( .A(B[0]), .B(A[0]), .Y(n2852) );
  XOR2X1 U2495 ( .A(n1660), .B(n147), .Y(SUM[50]) );
  INVX2 U2496 ( .A(n4698), .Y(n2911) );
  INVX2 U2497 ( .A(n4698), .Y(n3740) );
  INVX1 U2498 ( .A(n4652), .Y(n4738) );
  INVX8 U2499 ( .A(n4652), .Y(n4791) );
  INVX1 U2500 ( .A(n7), .Y(n2853) );
  INVX1 U2501 ( .A(n2107), .Y(n2854) );
  XOR2X1 U2502 ( .A(n2099), .B(n194), .Y(SUM[3]) );
  BUFX4 U2503 ( .A(n2900), .Y(n4698) );
  INVX1 U2504 ( .A(n4176), .Y(n2855) );
  INVX1 U2505 ( .A(n4477), .Y(n2856) );
  BUFX2 U2506 ( .A(n3526), .Y(n2857) );
  BUFX2 U2507 ( .A(n1750), .Y(n2858) );
  AND2X2 U2508 ( .A(n1780), .B(n1773), .Y(n2859) );
  OAI21X1 U2509 ( .A(n3465), .B(n3228), .C(n3151), .Y(n2860) );
  INVX1 U2510 ( .A(n2837), .Y(n4728) );
  INVX1 U2511 ( .A(n3398), .Y(n1966) );
  INVX1 U2512 ( .A(n4750), .Y(n4748) );
  INVX1 U2513 ( .A(n2951), .Y(n2181) );
  XOR2X1 U2514 ( .A(n2836), .B(n181), .Y(SUM[16]) );
  XNOR2X1 U2515 ( .A(n3740), .B(n165), .Y(SUM[32]) );
  INVX2 U2516 ( .A(n2898), .Y(n4643) );
  BUFX2 U2517 ( .A(n1643), .Y(n2861) );
  AND2X2 U2518 ( .A(n2949), .B(n406), .Y(n4782) );
  AND2X2 U2519 ( .A(n2048), .B(n2041), .Y(n2862) );
  INVX1 U2520 ( .A(n4652), .Y(n2863) );
  INVX1 U2521 ( .A(n4652), .Y(n2864) );
  INVX1 U2522 ( .A(n2910), .Y(n2865) );
  INVX1 U2523 ( .A(n4768), .Y(n2866) );
  INVX1 U2524 ( .A(n1840), .Y(n2867) );
  INVX1 U2525 ( .A(n4652), .Y(n2868) );
  INVX1 U2526 ( .A(n4652), .Y(n2869) );
  INVX1 U2527 ( .A(n3603), .Y(n2870) );
  INVX1 U2528 ( .A(n4176), .Y(n2871) );
  INVX1 U2529 ( .A(n1603), .Y(n2872) );
  INVX1 U2530 ( .A(n2003), .Y(n2873) );
  INVX1 U2531 ( .A(n4787), .Y(n2874) );
  INVX1 U2532 ( .A(n2874), .Y(n2875) );
  INVX1 U2533 ( .A(n4652), .Y(n2876) );
  INVX1 U2534 ( .A(n4694), .Y(n2877) );
  INVX1 U2535 ( .A(n1601), .Y(n2878) );
  INVX8 U2536 ( .A(n4787), .Y(n4793) );
  AND2X2 U2537 ( .A(n3728), .B(n2842), .Y(n2879) );
  INVX1 U2538 ( .A(n1477), .Y(n2880) );
  OAI21X1 U2539 ( .A(n4217), .B(n3503), .C(n3155), .Y(n2881) );
  INVX1 U2540 ( .A(n614), .Y(n2882) );
  INVX1 U2541 ( .A(n1164), .Y(n2883) );
  AND2X2 U2542 ( .A(n4714), .B(n1422), .Y(n2884) );
  INVX1 U2543 ( .A(n2884), .Y(n4316) );
  INVX1 U2544 ( .A(n4458), .Y(n2885) );
  INVX1 U2545 ( .A(n1256), .Y(n2886) );
  INVX4 U2546 ( .A(n3727), .Y(n1681) );
  INVX1 U2547 ( .A(n1972), .Y(n2887) );
  INVX8 U2548 ( .A(n4652), .Y(n2888) );
  INVX1 U2549 ( .A(n4652), .Y(n2889) );
  INVX1 U2550 ( .A(n1780), .Y(n2890) );
  INVX1 U2551 ( .A(n2890), .Y(n2891) );
  BUFX2 U2552 ( .A(n1401), .Y(n2892) );
  OAI21X1 U2553 ( .A(n3595), .B(n3534), .C(n3159), .Y(n2893) );
  INVX1 U2554 ( .A(n1160), .Y(n2894) );
  AND2X2 U2555 ( .A(n1160), .B(n1332), .Y(n2895) );
  INVX1 U2556 ( .A(n784), .Y(n2896) );
  OAI21X1 U2557 ( .A(n2866), .B(n3514), .C(n3288), .Y(n2897) );
  BUFX2 U2558 ( .A(n1764), .Y(n2898) );
  OAI21X1 U2559 ( .A(n3505), .B(n2894), .C(n3158), .Y(n2899) );
  OAI21X1 U2560 ( .A(n3465), .B(n3228), .C(n3151), .Y(n2900) );
  OR2X2 U2561 ( .A(n4792), .B(n3056), .Y(n1029) );
  XNOR2X1 U2562 ( .A(n1590), .B(n4007), .Y(SUM[56]) );
  AND2X2 U2563 ( .A(n3275), .B(n1506), .Y(n2901) );
  INVX2 U2564 ( .A(n3275), .Y(n1595) );
  OR2X2 U2565 ( .A(A[149]), .B(B[149]), .Y(n530) );
  INVX1 U2566 ( .A(n1338), .Y(n2902) );
  INVX1 U2567 ( .A(n1212), .Y(n2903) );
  AND2X2 U2568 ( .A(n964), .B(n744), .Y(n2904) );
  INVX1 U2569 ( .A(n3588), .Y(n2905) );
  INVX4 U2570 ( .A(n4651), .Y(n1682) );
  AND2X2 U2571 ( .A(n1805), .B(n1769), .Y(n2906) );
  BUFX2 U2572 ( .A(n748), .Y(n2907) );
  INVX1 U2573 ( .A(n1864), .Y(n2908) );
  INVX1 U2574 ( .A(n7), .Y(n2909) );
  INVX1 U2575 ( .A(n7), .Y(n2910) );
  AND2X2 U2576 ( .A(n1687), .B(n1725), .Y(n2912) );
  AND2X2 U2577 ( .A(n2850), .B(n888), .Y(n2913) );
  OR2X2 U2578 ( .A(n4792), .B(n3444), .Y(n875) );
  OR2X2 U2579 ( .A(n4792), .B(n3446), .Y(n858) );
  INVX8 U2580 ( .A(n2849), .Y(n4792) );
  OR2X2 U2581 ( .A(A[93]), .B(B[93]), .Y(n4166) );
  INVX1 U2582 ( .A(n4166), .Y(n2914) );
  AND2X2 U2583 ( .A(B[20]), .B(A[20]), .Y(n4211) );
  INVX1 U2584 ( .A(n4211), .Y(n2915) );
  AND2X2 U2585 ( .A(B[68]), .B(A[68]), .Y(n4212) );
  INVX1 U2586 ( .A(n4212), .Y(n2916) );
  AND2X2 U2587 ( .A(B[132]), .B(A[132]), .Y(n4214) );
  INVX1 U2588 ( .A(n4214), .Y(n2917) );
  AND2X2 U2589 ( .A(B[166]), .B(A[166]), .Y(n4215) );
  INVX1 U2590 ( .A(n4215), .Y(n2918) );
  AND2X2 U2591 ( .A(B[54]), .B(A[54]), .Y(n4221) );
  INVX1 U2592 ( .A(n4221), .Y(n2919) );
  AND2X2 U2593 ( .A(B[56]), .B(A[56]), .Y(n4222) );
  INVX1 U2594 ( .A(n4222), .Y(n2920) );
  AND2X2 U2595 ( .A(A[66]), .B(B[66]), .Y(n4223) );
  INVX1 U2596 ( .A(n4223), .Y(n2921) );
  AND2X2 U2597 ( .A(B[74]), .B(A[74]), .Y(n4226) );
  INVX1 U2598 ( .A(n4226), .Y(n2922) );
  AND2X2 U2599 ( .A(B[134]), .B(A[134]), .Y(n4229) );
  INVX1 U2600 ( .A(n4229), .Y(n2923) );
  AND2X2 U2601 ( .A(n2973), .B(n4242), .Y(n172) );
  INVX1 U2602 ( .A(n172), .Y(n2924) );
  OR2X2 U2603 ( .A(n3734), .B(n4703), .Y(n1630) );
  INVX1 U2604 ( .A(n1630), .Y(n2925) );
  OR2X2 U2605 ( .A(n3336), .B(n4721), .Y(n1608) );
  INVX1 U2606 ( .A(n1608), .Y(n2926) );
  OR2X2 U2607 ( .A(n1456), .B(n4446), .Y(n1447) );
  INVX1 U2608 ( .A(n1447), .Y(n2927) );
  AND2X2 U2609 ( .A(B[82]), .B(A[82]), .Y(n1310) );
  INVX1 U2610 ( .A(n1310), .Y(n2928) );
  OR2X2 U2611 ( .A(n1250), .B(n1230), .Y(n1228) );
  INVX1 U2612 ( .A(n1228), .Y(n2929) );
  OR2X2 U2613 ( .A(n1250), .B(n4772), .Y(n1204) );
  INVX1 U2614 ( .A(n1204), .Y(n2930) );
  AND2X2 U2615 ( .A(B[92]), .B(A[92]), .Y(n1198) );
  INVX1 U2616 ( .A(n1198), .Y(n2931) );
  OR2X2 U2617 ( .A(n1250), .B(n4301), .Y(n1182) );
  INVX1 U2618 ( .A(n1182), .Y(n2932) );
  OR2X2 U2619 ( .A(n4792), .B(n1088), .Y(n1086) );
  OR2X2 U2620 ( .A(n4792), .B(n4304), .Y(n1077) );
  INVX1 U2621 ( .A(n1077), .Y(n2933) );
  OR2X2 U2622 ( .A(n4792), .B(n3066), .Y(n979) );
  INVX1 U2623 ( .A(n979), .Y(n2934) );
  OR2X2 U2624 ( .A(n944), .B(n4399), .Y(n933) );
  INVX1 U2625 ( .A(n933), .Y(n2935) );
  OR2X2 U2626 ( .A(n4792), .B(n3437), .Y(n929) );
  INVX1 U2627 ( .A(n929), .Y(n2936) );
  OR2X2 U2628 ( .A(n4792), .B(n3439), .Y(n912) );
  INVX1 U2629 ( .A(n912), .Y(n2937) );
  OR2X2 U2630 ( .A(n4319), .B(n4377), .Y(n905) );
  INVX1 U2631 ( .A(n905), .Y(n2938) );
  OR2X2 U2632 ( .A(n4792), .B(n3441), .Y(n901) );
  INVX1 U2633 ( .A(n901), .Y(n2939) );
  OR2X2 U2634 ( .A(n4792), .B(n3450), .Y(n830) );
  INVX1 U2635 ( .A(n830), .Y(n2940) );
  OR2X2 U2636 ( .A(n4792), .B(n3452), .Y(n817) );
  INVX1 U2637 ( .A(n817), .Y(n2941) );
  AND2X2 U2638 ( .A(B[146]), .B(A[146]), .Y(n562) );
  INVX1 U2639 ( .A(n562), .Y(n2942) );
  OR2X2 U2640 ( .A(n3738), .B(n526), .Y(n524) );
  INVX1 U2641 ( .A(n524), .Y(n2943) );
  OR2X2 U2642 ( .A(n3118), .B(n4366), .Y(n445) );
  INVX1 U2643 ( .A(n445), .Y(n2944) );
  OR2X2 U2644 ( .A(n3178), .B(n3599), .Y(n414) );
  INVX1 U2645 ( .A(n414), .Y(n2945) );
  OR2X2 U2646 ( .A(n408), .B(n4615), .Y(n399) );
  INVX1 U2647 ( .A(n399), .Y(n2946) );
  OR2X2 U2648 ( .A(n3464), .B(n352), .Y(n348) );
  INVX1 U2649 ( .A(n348), .Y(n2947) );
  OR2X2 U2650 ( .A(n324), .B(n3753), .Y(n304) );
  INVX1 U2651 ( .A(n304), .Y(n2948) );
  OR2X2 U2652 ( .A(n3364), .B(n4313), .Y(n205) );
  INVX1 U2653 ( .A(n205), .Y(n2949) );
  OR2X2 U2654 ( .A(A[49]), .B(B[49]), .Y(n3886) );
  OR2X2 U2655 ( .A(A[28]), .B(B[28]), .Y(n4148) );
  AND2X2 U2656 ( .A(n4288), .B(n406), .Y(n4163) );
  INVX1 U2657 ( .A(n4163), .Y(n2950) );
  OR2X2 U2658 ( .A(A[26]), .B(B[26]), .Y(n4168) );
  OR2X2 U2659 ( .A(A[44]), .B(B[44]), .Y(n4170) );
  OR2X2 U2660 ( .A(A[54]), .B(B[54]), .Y(n4173) );
  OR2X2 U2661 ( .A(A[72]), .B(B[72]), .Y(n4175) );
  OR2X2 U2662 ( .A(A[77]), .B(B[77]), .Y(n4176) );
  OR2X2 U2663 ( .A(A[91]), .B(B[91]), .Y(n4178) );
  OR2X2 U2664 ( .A(A[101]), .B(B[101]), .Y(n4180) );
  OR2X2 U2665 ( .A(A[102]), .B(B[102]), .Y(n4181) );
  OR2X2 U2666 ( .A(A[106]), .B(B[106]), .Y(n4182) );
  INVX1 U2667 ( .A(n4182), .Y(n2951) );
  OR2X2 U2668 ( .A(A[107]), .B(B[107]), .Y(n4183) );
  INVX1 U2669 ( .A(n4183), .Y(n2952) );
  OR2X2 U2670 ( .A(A[110]), .B(B[110]), .Y(n4184) );
  OR2X2 U2671 ( .A(A[119]), .B(B[119]), .Y(n4185) );
  OR2X2 U2672 ( .A(A[25]), .B(B[25]), .Y(n4242) );
  OR2X2 U2673 ( .A(A[97]), .B(B[97]), .Y(n4247) );
  OR2X2 U2674 ( .A(A[133]), .B(B[133]), .Y(n4250) );
  OR2X2 U2675 ( .A(A[157]), .B(B[157]), .Y(n4251) );
  INVX1 U2676 ( .A(n4251), .Y(n2953) );
  OR2X2 U2677 ( .A(A[173]), .B(B[173]), .Y(n4252) );
  INVX1 U2678 ( .A(n4252), .Y(n2954) );
  AND2X2 U2679 ( .A(B[94]), .B(A[94]), .Y(n4331) );
  INVX1 U2680 ( .A(n4331), .Y(n2955) );
  AND2X2 U2681 ( .A(B[100]), .B(A[100]), .Y(n4345) );
  OR2X2 U2682 ( .A(A[73]), .B(B[73]), .Y(n4458) );
  OR2X2 U2683 ( .A(A[53]), .B(B[53]), .Y(n4480) );
  OR2X2 U2684 ( .A(A[109]), .B(B[109]), .Y(n4497) );
  OR2X2 U2685 ( .A(A[114]), .B(B[114]), .Y(n4704) );
  AND2X2 U2686 ( .A(n3323), .B(n3890), .Y(n4705) );
  OR2X2 U2687 ( .A(A[76]), .B(B[76]), .Y(n4758) );
  OR2X2 U2688 ( .A(A[33]), .B(B[33]), .Y(n4768) );
  AND2X2 U2689 ( .A(B[1]), .B(A[1]), .Y(n2105) );
  INVX1 U2690 ( .A(n2105), .Y(n2956) );
  AND2X2 U2691 ( .A(B[3]), .B(A[3]), .Y(n2098) );
  INVX1 U2692 ( .A(n2098), .Y(n2957) );
  AND2X2 U2693 ( .A(B[5]), .B(A[5]), .Y(n2087) );
  INVX1 U2694 ( .A(n2087), .Y(n2958) );
  AND2X2 U2695 ( .A(B[6]), .B(A[6]), .Y(n2078) );
  INVX1 U2696 ( .A(n2078), .Y(n2959) );
  AND2X2 U2697 ( .A(B[7]), .B(A[7]), .Y(n2071) );
  INVX1 U2698 ( .A(n2071), .Y(n2960) );
  OR2X2 U2699 ( .A(A[8]), .B(B[8]), .Y(n2062) );
  INVX1 U2700 ( .A(n2062), .Y(n2961) );
  AND2X2 U2701 ( .A(B[9]), .B(A[9]), .Y(n2060) );
  INVX1 U2702 ( .A(n2060), .Y(n2962) );
  AND2X2 U2703 ( .A(B[11]), .B(A[11]), .Y(n2042) );
  INVX1 U2704 ( .A(n2042), .Y(n2963) );
  OR2X2 U2705 ( .A(A[13]), .B(B[13]), .Y(n2023) );
  OR2X2 U2706 ( .A(A[15]), .B(B[15]), .Y(n2003) );
  INVX1 U2707 ( .A(n2003), .Y(n2964) );
  OR2X2 U2708 ( .A(n3330), .B(n3589), .Y(n1997) );
  AND2X2 U2709 ( .A(B[17]), .B(A[17]), .Y(n1989) );
  INVX1 U2710 ( .A(n1989), .Y(n2965) );
  AND2X2 U2711 ( .A(B[18]), .B(A[18]), .Y(n1980) );
  INVX1 U2712 ( .A(n1980), .Y(n2966) );
  AND2X2 U2713 ( .A(B[19]), .B(A[19]), .Y(n1973) );
  INVX1 U2714 ( .A(n1973), .Y(n2967) );
  OR2X2 U2715 ( .A(A[19]), .B(B[19]), .Y(n1972) );
  INVX1 U2716 ( .A(n1972), .Y(n2968) );
  OR2X2 U2717 ( .A(n2887), .B(n4779), .Y(n1970) );
  AND2X2 U2718 ( .A(B[21]), .B(A[21]), .Y(n1953) );
  INVX1 U2719 ( .A(n1953), .Y(n2969) );
  AND2X2 U2720 ( .A(B[22]), .B(A[22]), .Y(n1942) );
  INVX1 U2721 ( .A(n1942), .Y(n2970) );
  OR2X2 U2722 ( .A(A[23]), .B(B[23]), .Y(n1934) );
  INVX1 U2723 ( .A(n1934), .Y(n2971) );
  OR2X2 U2724 ( .A(A[24]), .B(B[24]), .Y(n1919) );
  OR2X1 U2725 ( .A(n1926), .B(n4661), .Y(n1917) );
  INVX1 U2726 ( .A(n1917), .Y(n2972) );
  AND2X2 U2727 ( .A(B[25]), .B(A[25]), .Y(n1915) );
  INVX1 U2728 ( .A(n1915), .Y(n2973) );
  OR2X2 U2729 ( .A(n1926), .B(n1906), .Y(n1904) );
  INVX1 U2730 ( .A(n1904), .Y(n2974) );
  AND2X2 U2731 ( .A(B[26]), .B(A[26]), .Y(n1902) );
  INVX1 U2732 ( .A(n1902), .Y(n2975) );
  OR2X2 U2733 ( .A(n1926), .B(n4292), .Y(n1895) );
  INVX1 U2734 ( .A(n1895), .Y(n2976) );
  AND2X2 U2735 ( .A(B[27]), .B(A[27]), .Y(n1893) );
  INVX1 U2736 ( .A(n1893), .Y(n2977) );
  OR2X2 U2737 ( .A(n3174), .B(n3405), .Y(n1890) );
  INVX1 U2738 ( .A(n1890), .Y(n2978) );
  OR2X1 U2739 ( .A(n1926), .B(n4752), .Y(n1882) );
  INVX1 U2740 ( .A(n1882), .Y(n2979) );
  OR2X1 U2741 ( .A(n1926), .B(n4293), .Y(n1873) );
  INVX1 U2742 ( .A(n1873), .Y(n2980) );
  AND2X2 U2743 ( .A(B[29]), .B(A[29]), .Y(n1871) );
  INVX1 U2744 ( .A(n1871), .Y(n2981) );
  OR2X2 U2745 ( .A(A[29]), .B(B[29]), .Y(n1870) );
  INVX1 U2746 ( .A(n1870), .Y(n2982) );
  OR2X2 U2747 ( .A(n3866), .B(n2982), .Y(n1864) );
  INVX1 U2748 ( .A(n1864), .Y(n2983) );
  OR2X1 U2749 ( .A(n1926), .B(n4294), .Y(n1860) );
  INVX1 U2750 ( .A(n1860), .Y(n2984) );
  AND2X2 U2751 ( .A(B[30]), .B(A[30]), .Y(n1858) );
  INVX1 U2752 ( .A(n1858), .Y(n2985) );
  OR2X1 U2753 ( .A(n1926), .B(n4295), .Y(n1849) );
  INVX1 U2754 ( .A(n1849), .Y(n2986) );
  AND2X2 U2755 ( .A(B[31]), .B(A[31]), .Y(n1847) );
  INVX1 U2756 ( .A(n1847), .Y(n2987) );
  OR2X2 U2757 ( .A(A[31]), .B(B[31]), .Y(n1846) );
  OR2X2 U2758 ( .A(n3333), .B(n3415), .Y(n1840) );
  OR2X2 U2759 ( .A(n2866), .B(n3417), .Y(n1825) );
  INVX1 U2760 ( .A(n1825), .Y(n2988) );
  AND2X2 U2761 ( .A(B[35]), .B(A[35]), .Y(n1814) );
  INVX1 U2762 ( .A(n1814), .Y(n2989) );
  AND2X2 U2763 ( .A(B[36]), .B(A[36]), .Y(n1799) );
  INVX1 U2764 ( .A(n1799), .Y(n2990) );
  OR2X2 U2765 ( .A(A[37]), .B(B[37]), .Y(n1791) );
  AND2X2 U2766 ( .A(B[38]), .B(A[38]), .Y(n1781) );
  INVX1 U2767 ( .A(n1781), .Y(n2991) );
  AND2X2 U2768 ( .A(B[39]), .B(A[39]), .Y(n1774) );
  INVX1 U2769 ( .A(n1774), .Y(n2992) );
  AND2X2 U2770 ( .A(n2859), .B(n3297), .Y(n1769) );
  INVX1 U2771 ( .A(n1769), .Y(n2993) );
  OR2X2 U2772 ( .A(A[40]), .B(B[40]), .Y(n1758) );
  AND2X2 U2773 ( .A(A[41]), .B(B[41]), .Y(n1752) );
  INVX1 U2774 ( .A(n1752), .Y(n2994) );
  OR2X2 U2775 ( .A(A[42]), .B(B[42]), .Y(n1740) );
  AND2X2 U2776 ( .A(B[43]), .B(A[43]), .Y(n1734) );
  INVX1 U2777 ( .A(n1734), .Y(n2995) );
  OR2X2 U2778 ( .A(A[43]), .B(B[43]), .Y(n1733) );
  INVX1 U2779 ( .A(n1733), .Y(n2996) );
  AND2X2 U2780 ( .A(B[44]), .B(A[44]), .Y(n1719) );
  INVX1 U2781 ( .A(n1719), .Y(n2997) );
  AND2X2 U2782 ( .A(B[45]), .B(A[45]), .Y(n1712) );
  INVX1 U2783 ( .A(n1712), .Y(n2998) );
  AND2X2 U2784 ( .A(B[46]), .B(A[46]), .Y(n1699) );
  INVX1 U2785 ( .A(n1699), .Y(n2999) );
  AND2X2 U2786 ( .A(B[47]), .B(A[47]), .Y(n1692) );
  INVX1 U2787 ( .A(n1692), .Y(n3000) );
  OR2X2 U2788 ( .A(A[48]), .B(B[48]), .Y(n1676) );
  AND2X2 U2789 ( .A(B[49]), .B(A[49]), .Y(n1670) );
  INVX1 U2790 ( .A(n1670), .Y(n3001) );
  OR2X2 U2791 ( .A(n3170), .B(n3870), .Y(n1663) );
  OR2X2 U2792 ( .A(A[50]), .B(B[50]), .Y(n1656) );
  AND2X2 U2793 ( .A(B[51]), .B(A[51]), .Y(n1650) );
  INVX1 U2794 ( .A(n1650), .Y(n3002) );
  OR2X2 U2795 ( .A(A[51]), .B(B[51]), .Y(n1649) );
  OR2X2 U2796 ( .A(n3171), .B(n4449), .Y(n1647) );
  AND2X2 U2797 ( .A(B[52]), .B(A[52]), .Y(n1635) );
  OR2X2 U2798 ( .A(A[52]), .B(B[52]), .Y(n1632) );
  AND2X2 U2799 ( .A(B[53]), .B(A[53]), .Y(n1626) );
  INVX1 U2800 ( .A(n1626), .Y(n3003) );
  OR2X2 U2801 ( .A(n3871), .B(n4172), .Y(n1621) );
  AND2X2 U2802 ( .A(B[55]), .B(A[55]), .Y(n1604) );
  INVX1 U2803 ( .A(n1604), .Y(n3004) );
  OR2X2 U2804 ( .A(A[55]), .B(B[55]), .Y(n1603) );
  INVX1 U2805 ( .A(n1603), .Y(n3005) );
  OR2X2 U2806 ( .A(n3901), .B(n2872), .Y(n1601) );
  INVX1 U2807 ( .A(n1601), .Y(n3006) );
  OR2X2 U2808 ( .A(n1595), .B(n4711), .Y(n1584) );
  INVX1 U2809 ( .A(n1584), .Y(n3007) );
  AND2X2 U2810 ( .A(B[57]), .B(A[57]), .Y(n1580) );
  INVX1 U2811 ( .A(n1580), .Y(n3008) );
  OR2X2 U2812 ( .A(A[57]), .B(B[57]), .Y(n1579) );
  OR2X2 U2813 ( .A(n1595), .B(n1571), .Y(n1569) );
  INVX1 U2814 ( .A(n1569), .Y(n3009) );
  OR2X1 U2815 ( .A(n1595), .B(n4297), .Y(n1558) );
  INVX1 U2816 ( .A(n1558), .Y(n3010) );
  AND2X2 U2817 ( .A(B[59]), .B(A[59]), .Y(n1554) );
  INVX1 U2818 ( .A(n1554), .Y(n3011) );
  OR2X2 U2819 ( .A(A[59]), .B(B[59]), .Y(n1553) );
  OR2X2 U2820 ( .A(n1595), .B(n4742), .Y(n1543) );
  INVX1 U2821 ( .A(n1543), .Y(n3012) );
  OR2X1 U2822 ( .A(n1595), .B(n4298), .Y(n1532) );
  INVX1 U2823 ( .A(n1532), .Y(n3013) );
  AND2X2 U2824 ( .A(B[61]), .B(A[61]), .Y(n1528) );
  INVX1 U2825 ( .A(n1528), .Y(n3014) );
  OR2X2 U2826 ( .A(A[61]), .B(B[61]), .Y(n1527) );
  INVX1 U2827 ( .A(n1527), .Y(n3015) );
  OR2X2 U2828 ( .A(n1595), .B(n4299), .Y(n1517) );
  INVX1 U2829 ( .A(n1517), .Y(n3016) );
  AND2X2 U2830 ( .A(B[62]), .B(A[62]), .Y(n1513) );
  OR2X2 U2831 ( .A(A[62]), .B(B[62]), .Y(n1510) );
  INVX1 U2832 ( .A(n1510), .Y(n3017) );
  AND2X2 U2833 ( .A(B[63]), .B(A[63]), .Y(n1500) );
  INVX1 U2834 ( .A(n1500), .Y(n3018) );
  OR2X2 U2835 ( .A(A[63]), .B(B[63]), .Y(n1499) );
  OR2X2 U2836 ( .A(n3339), .B(n3427), .Y(n1493) );
  OR2X2 U2837 ( .A(n3574), .B(n3726), .Y(n1489) );
  AND2X2 U2838 ( .A(B[65]), .B(A[65]), .Y(n1481) );
  INVX1 U2839 ( .A(n1481), .Y(n3019) );
  AND2X2 U2840 ( .A(B[67]), .B(A[67]), .Y(n1465) );
  INVX1 U2841 ( .A(n1465), .Y(n3020) );
  OR2X2 U2842 ( .A(A[69]), .B(B[69]), .Y(n1444) );
  OR2X2 U2843 ( .A(A[71]), .B(B[71]), .Y(n1426) );
  OR2X2 U2844 ( .A(n3754), .B(n4456), .Y(n1424) );
  INVX1 U2845 ( .A(n1424), .Y(n3021) );
  AND2X2 U2846 ( .A(n3021), .B(n3299), .Y(n1422) );
  AND2X2 U2847 ( .A(B[73]), .B(A[73]), .Y(n1403) );
  INVX1 U2848 ( .A(n1403), .Y(n3022) );
  OR2X2 U2849 ( .A(n3902), .B(n2885), .Y(n1398) );
  OR2X2 U2850 ( .A(A[74]), .B(B[74]), .Y(n1389) );
  INVX1 U2851 ( .A(n1389), .Y(n3023) );
  AND2X2 U2852 ( .A(B[75]), .B(A[75]), .Y(n1385) );
  INVX1 U2853 ( .A(n1385), .Y(n3024) );
  OR2X2 U2854 ( .A(A[75]), .B(B[75]), .Y(n1384) );
  OR2X2 U2855 ( .A(n3023), .B(n4459), .Y(n1382) );
  OR2X2 U2856 ( .A(n4316), .B(n3325), .Y(n1372) );
  INVX1 U2857 ( .A(n1372), .Y(n3025) );
  AND2X2 U2858 ( .A(B[77]), .B(A[77]), .Y(n1363) );
  INVX1 U2859 ( .A(n1363), .Y(n3026) );
  AND2X2 U2860 ( .A(B[78]), .B(A[78]), .Y(n1352) );
  INVX1 U2861 ( .A(n1352), .Y(n3027) );
  OR2X2 U2862 ( .A(n1340), .B(n3324), .Y(n1338) );
  OR2X2 U2863 ( .A(A[81]), .B(B[81]), .Y(n1320) );
  OR2X2 U2864 ( .A(n3175), .B(n3401), .Y(n1300) );
  INVX1 U2865 ( .A(n1300), .Y(n3028) );
  AND2X2 U2866 ( .A(n3028), .B(n3289), .Y(n1294) );
  AND2X2 U2867 ( .A(n1292), .B(n2848), .Y(n1290) );
  INVX1 U2868 ( .A(n1290), .Y(n3029) );
  AND2X2 U2869 ( .A(B[84]), .B(A[84]), .Y(n1286) );
  INVX1 U2870 ( .A(n1286), .Y(n3030) );
  OR2X2 U2871 ( .A(A[87]), .B(B[87]), .Y(n1258) );
  INVX1 U2872 ( .A(n1258), .Y(n3031) );
  OR2X2 U2873 ( .A(n4177), .B(n3201), .Y(n1256) );
  INVX1 U2874 ( .A(n1256), .Y(n3032) );
  OR2X2 U2875 ( .A(A[89]), .B(B[89]), .Y(n1234) );
  AND2X2 U2876 ( .A(B[90]), .B(A[90]), .Y(n1222) );
  INVX1 U2877 ( .A(n1222), .Y(n3033) );
  OR2X2 U2878 ( .A(A[90]), .B(B[90]), .Y(n1219) );
  OR2X2 U2879 ( .A(n3875), .B(n4729), .Y(n1217) );
  INVX1 U2880 ( .A(n1217), .Y(n3034) );
  AND2X2 U2881 ( .A(B[91]), .B(A[91]), .Y(n1215) );
  INVX1 U2882 ( .A(n1215), .Y(n3035) );
  OR2X2 U2883 ( .A(n3910), .B(n4154), .Y(n1212) );
  INVX1 U2884 ( .A(n1212), .Y(n3036) );
  OR2X2 U2885 ( .A(n3877), .B(n4438), .Y(n1193) );
  INVX1 U2886 ( .A(n1193), .Y(n3037) );
  OR2X2 U2887 ( .A(n4155), .B(n4734), .Y(n1171) );
  INVX1 U2888 ( .A(n1171), .Y(n3038) );
  AND2X2 U2889 ( .A(B[95]), .B(A[95]), .Y(n1169) );
  INVX1 U2890 ( .A(n1169), .Y(n3039) );
  AND2X2 U2891 ( .A(n3311), .B(n3291), .Y(n1164) );
  INVX1 U2892 ( .A(n1164), .Y(n3040) );
  AND2X2 U2893 ( .A(n3301), .B(n3313), .Y(n1160) );
  OR2X2 U2894 ( .A(A[96]), .B(B[96]), .Y(n1149) );
  OR2X2 U2895 ( .A(n4792), .B(n4601), .Y(n1147) );
  INVX1 U2896 ( .A(n1147), .Y(n3041) );
  AND2X2 U2897 ( .A(B[97]), .B(A[97]), .Y(n1145) );
  INVX1 U2898 ( .A(n1145), .Y(n3042) );
  OR2X2 U2899 ( .A(A[98]), .B(B[98]), .Y(n1131) );
  INVX1 U2900 ( .A(n1131), .Y(n3043) );
  OR2X2 U2901 ( .A(n4792), .B(n4302), .Y(n1125) );
  INVX1 U2902 ( .A(n1125), .Y(n3044) );
  AND2X2 U2903 ( .A(B[99]), .B(A[99]), .Y(n1123) );
  INVX1 U2904 ( .A(n1123), .Y(n3045) );
  OR2X2 U2905 ( .A(A[99]), .B(B[99]), .Y(n1122) );
  INVX1 U2906 ( .A(n1122), .Y(n3046) );
  OR2X2 U2907 ( .A(n4723), .B(n4792), .Y(n1108) );
  INVX1 U2908 ( .A(n1108), .Y(n3047) );
  OR2X2 U2909 ( .A(n4792), .B(n4303), .Y(n1099) );
  INVX1 U2910 ( .A(n1099), .Y(n3048) );
  AND2X2 U2911 ( .A(B[101]), .B(A[101]), .Y(n1097) );
  INVX1 U2912 ( .A(n1097), .Y(n3049) );
  AND2X2 U2913 ( .A(B[103]), .B(A[103]), .Y(n1075) );
  INVX1 U2914 ( .A(n1075), .Y(n3050) );
  OR2X2 U2915 ( .A(n3176), .B(n3433), .Y(n1072) );
  INVX1 U2916 ( .A(n1072), .Y(n3051) );
  OR2X2 U2917 ( .A(n3735), .B(n3596), .Y(n1064) );
  INVX1 U2918 ( .A(n1064), .Y(n3052) );
  OR2X2 U2919 ( .A(n4792), .B(n1064), .Y(n1060) );
  INVX1 U2920 ( .A(n1060), .Y(n3053) );
  OR2X2 U2921 ( .A(n4792), .B(n4305), .Y(n1051) );
  INVX1 U2922 ( .A(n1051), .Y(n3054) );
  OR2X2 U2923 ( .A(A[105]), .B(B[105]), .Y(n1048) );
  OR2X2 U2924 ( .A(n4792), .B(n1040), .Y(n1038) );
  INVX1 U2925 ( .A(n1038), .Y(n3055) );
  AND2X2 U2926 ( .A(B[106]), .B(A[106]), .Y(n1036) );
  AND2X2 U2927 ( .A(n2181), .B(n4137), .Y(n1031) );
  INVX1 U2928 ( .A(n1031), .Y(n3056) );
  INVX1 U2929 ( .A(n1029), .Y(n3057) );
  AND2X2 U2930 ( .A(B[107]), .B(A[107]), .Y(n1027) );
  INVX1 U2931 ( .A(n1027), .Y(n3058) );
  OR2X2 U2932 ( .A(n2951), .B(n2952), .Y(n1024) );
  AND2X2 U2933 ( .A(n4283), .B(n3303), .Y(n1018) );
  OR2X1 U2934 ( .A(n4792), .B(n1014), .Y(n1012) );
  INVX1 U2935 ( .A(n1012), .Y(n3059) );
  AND2X2 U2936 ( .A(B[108]), .B(A[108]), .Y(n1010) );
  OR2X2 U2937 ( .A(A[108]), .B(B[108]), .Y(n1009) );
  INVX1 U2938 ( .A(n1009), .Y(n3060) );
  AND2X2 U2939 ( .A(n1009), .B(n3304), .Y(n1005) );
  INVX1 U2940 ( .A(n1005), .Y(n3061) );
  OR2X1 U2941 ( .A(n4792), .B(n3061), .Y(n1003) );
  INVX1 U2942 ( .A(n1003), .Y(n3062) );
  AND2X2 U2943 ( .A(B[109]), .B(A[109]), .Y(n1001) );
  INVX1 U2944 ( .A(n1001), .Y(n3063) );
  OR2X2 U2945 ( .A(n3060), .B(n3911), .Y(n996) );
  INVX1 U2946 ( .A(n996), .Y(n3064) );
  OR2X2 U2947 ( .A(n4792), .B(n990), .Y(n988) );
  INVX1 U2948 ( .A(n988), .Y(n3065) );
  AND2X2 U2949 ( .A(n4184), .B(n3306), .Y(n981) );
  INVX1 U2950 ( .A(n981), .Y(n3066) );
  AND2X2 U2951 ( .A(B[111]), .B(A[111]), .Y(n977) );
  INVX1 U2952 ( .A(n977), .Y(n3067) );
  OR2X2 U2953 ( .A(n3344), .B(n3202), .Y(n974) );
  INVX1 U2954 ( .A(n974), .Y(n3068) );
  OR2X2 U2955 ( .A(n3326), .B(n4792), .Y(n962) );
  INVX1 U2956 ( .A(n962), .Y(n3069) );
  OR2X2 U2957 ( .A(A[112]), .B(B[112]), .Y(n959) );
  AND2X2 U2958 ( .A(n959), .B(n4689), .Y(n955) );
  INVX1 U2959 ( .A(n955), .Y(n3070) );
  OR2X2 U2960 ( .A(n4792), .B(n3070), .Y(n953) );
  INVX1 U2961 ( .A(n953), .Y(n3071) );
  AND2X2 U2962 ( .A(B[113]), .B(A[113]), .Y(n951) );
  INVX1 U2963 ( .A(n951), .Y(n3072) );
  OR2X2 U2964 ( .A(n3172), .B(n3436), .Y(n944) );
  AND2X2 U2965 ( .A(n4660), .B(n2879), .Y(n942) );
  INVX1 U2966 ( .A(n942), .Y(n3073) );
  OR2X2 U2967 ( .A(n4792), .B(n3073), .Y(n940) );
  INVX1 U2968 ( .A(n940), .Y(n3074) );
  AND2X2 U2969 ( .A(B[114]), .B(A[114]), .Y(n938) );
  AND2X2 U2970 ( .A(B[115]), .B(A[115]), .Y(n927) );
  INVX1 U2971 ( .A(n927), .Y(n3075) );
  OR2X2 U2972 ( .A(A[115]), .B(B[115]), .Y(n926) );
  AND2X2 U2973 ( .A(n3317), .B(n3874), .Y(n918) );
  AND2X2 U2974 ( .A(B[117]), .B(A[117]), .Y(n899) );
  INVX1 U2975 ( .A(n899), .Y(n3076) );
  OR2X2 U2976 ( .A(A[117]), .B(B[117]), .Y(n898) );
  OR2X2 U2977 ( .A(n4498), .B(n3912), .Y(n894) );
  INVX1 U2978 ( .A(n894), .Y(n3077) );
  OR2X2 U2979 ( .A(n3346), .B(n4389), .Y(n879) );
  INVX1 U2980 ( .A(n879), .Y(n3078) );
  AND2X2 U2981 ( .A(B[119]), .B(A[119]), .Y(n873) );
  INVX1 U2982 ( .A(n873), .Y(n3079) );
  OR2X2 U2983 ( .A(n3903), .B(n3868), .Y(n870) );
  INVX1 U2984 ( .A(n870), .Y(n3080) );
  AND2X2 U2985 ( .A(n3080), .B(n3077), .Y(n868) );
  INVX1 U2986 ( .A(n868), .Y(n3081) );
  OR2X2 U2987 ( .A(A[120]), .B(B[120]), .Y(n853) );
  OR2X2 U2988 ( .A(n4792), .B(n3449), .Y(n847) );
  INVX1 U2989 ( .A(n847), .Y(n3082) );
  AND2X2 U2990 ( .A(B[121]), .B(A[121]), .Y(n845) );
  INVX1 U2991 ( .A(n845), .Y(n3083) );
  OR2X2 U2992 ( .A(A[121]), .B(B[121]), .Y(n844) );
  AND2X2 U2993 ( .A(B[122]), .B(A[122]), .Y(n828) );
  OR2X2 U2994 ( .A(A[122]), .B(B[122]), .Y(n827) );
  AND2X2 U2995 ( .A(B[123]), .B(A[123]), .Y(n815) );
  INVX1 U2996 ( .A(n815), .Y(n3084) );
  OR2X2 U2997 ( .A(A[123]), .B(B[123]), .Y(n814) );
  OR2X2 U2998 ( .A(n4792), .B(n3455), .Y(n800) );
  INVX1 U2999 ( .A(n800), .Y(n3085) );
  OR2X2 U3000 ( .A(n4792), .B(n3457), .Y(n787) );
  INVX1 U3001 ( .A(n787), .Y(n3086) );
  AND2X2 U3002 ( .A(B[125]), .B(A[125]), .Y(n785) );
  INVX1 U3003 ( .A(n785), .Y(n3087) );
  OR2X2 U3004 ( .A(A[125]), .B(B[125]), .Y(n784) );
  OR2X2 U3005 ( .A(n4503), .B(n3234), .Y(n778) );
  OR2X2 U3006 ( .A(n4792), .B(n3459), .Y(n770) );
  INVX1 U3007 ( .A(n770), .Y(n3088) );
  OR2X2 U3008 ( .A(n4792), .B(n3461), .Y(n755) );
  INVX1 U3009 ( .A(n755), .Y(n3089) );
  AND2X2 U3010 ( .A(B[127]), .B(A[127]), .Y(n753) );
  INVX1 U3011 ( .A(n753), .Y(n3090) );
  OR2X2 U3012 ( .A(A[127]), .B(B[127]), .Y(n752) );
  INVX1 U3013 ( .A(n752), .Y(n3091) );
  OR2X2 U3014 ( .A(n3904), .B(n3091), .Y(n750) );
  OR2X2 U3015 ( .A(n3347), .B(n3402), .Y(n746) );
  INVX1 U3016 ( .A(n746), .Y(n3092) );
  OR2X2 U3017 ( .A(A[128]), .B(B[128]), .Y(n737) );
  OR2X2 U3018 ( .A(A[129]), .B(B[129]), .Y(n732) );
  AND2X2 U3019 ( .A(B[131]), .B(A[131]), .Y(n717) );
  INVX1 U3020 ( .A(n717), .Y(n3093) );
  OR2X2 U3021 ( .A(A[131]), .B(B[131]), .Y(n716) );
  INVX1 U3022 ( .A(n716), .Y(n3094) );
  AND2X2 U3023 ( .A(n3320), .B(n3307), .Y(n708) );
  AND2X2 U3024 ( .A(B[133]), .B(A[133]), .Y(n697) );
  INVX1 U3025 ( .A(n697), .Y(n3095) );
  OR2X2 U3026 ( .A(n4506), .B(n3913), .Y(n692) );
  AND2X2 U3027 ( .A(B[135]), .B(A[135]), .Y(n679) );
  INVX1 U3028 ( .A(n679), .Y(n3096) );
  OR2X2 U3029 ( .A(A[135]), .B(B[135]), .Y(n678) );
  INVX1 U3030 ( .A(n678), .Y(n3097) );
  OR2X2 U3031 ( .A(n3177), .B(n3097), .Y(n676) );
  INVX1 U3032 ( .A(n676), .Y(n3098) );
  OR2X2 U3033 ( .A(n4320), .B(n3597), .Y(n668) );
  AND2X2 U3034 ( .A(B[137]), .B(A[137]), .Y(n655) );
  INVX1 U3035 ( .A(n655), .Y(n3099) );
  OR2X2 U3036 ( .A(A[137]), .B(B[137]), .Y(n654) );
  OR2X2 U3037 ( .A(n4466), .B(n3914), .Y(n650) );
  AND2X2 U3038 ( .A(B[139]), .B(A[139]), .Y(n637) );
  INVX1 U3039 ( .A(n637), .Y(n3100) );
  OR2X2 U3040 ( .A(A[139]), .B(B[139]), .Y(n636) );
  INVX1 U3041 ( .A(n636), .Y(n3101) );
  OR2X2 U3042 ( .A(n3101), .B(n3869), .Y(n634) );
  INVX1 U3043 ( .A(n634), .Y(n3102) );
  AND2X2 U3044 ( .A(n3102), .B(n4541), .Y(n630) );
  INVX1 U3045 ( .A(n630), .Y(n3103) );
  AND2X2 U3046 ( .A(B[141]), .B(A[141]), .Y(n615) );
  INVX1 U3047 ( .A(n615), .Y(n3104) );
  OR2X2 U3048 ( .A(A[141]), .B(B[141]), .Y(n614) );
  OR2X2 U3049 ( .A(n4467), .B(n3915), .Y(n610) );
  INVX1 U3050 ( .A(n610), .Y(n3105) );
  AND2X2 U3051 ( .A(B[143]), .B(A[143]), .Y(n597) );
  INVX1 U3052 ( .A(n597), .Y(n3106) );
  OR2X2 U3053 ( .A(A[143]), .B(B[143]), .Y(n596) );
  INVX1 U3054 ( .A(n596), .Y(n3107) );
  OR2X2 U3055 ( .A(n3107), .B(n3916), .Y(n594) );
  INVX1 U3056 ( .A(n594), .Y(n3108) );
  AND2X2 U3057 ( .A(n3108), .B(n3105), .Y(n592) );
  INVX1 U3058 ( .A(n592), .Y(n3109) );
  OR2X2 U3059 ( .A(n3103), .B(n3109), .Y(n590) );
  INVX1 U3060 ( .A(n590), .Y(n3110) );
  OR2X2 U3061 ( .A(A[144]), .B(B[144]), .Y(n577) );
  OR2X2 U3062 ( .A(A[145]), .B(B[145]), .Y(n572) );
  OR2X2 U3063 ( .A(n4604), .B(n4187), .Y(n568) );
  INVX1 U3064 ( .A(n568), .Y(n3111) );
  OR2X2 U3065 ( .A(A[148]), .B(B[148]), .Y(n535) );
  AND2X2 U3066 ( .A(B[150]), .B(A[150]), .Y(n518) );
  INVX1 U3067 ( .A(n518), .Y(n3112) );
  AND2X2 U3068 ( .A(n3321), .B(n3309), .Y(n506) );
  INVX1 U3069 ( .A(n506), .Y(n3113) );
  OR2X2 U3070 ( .A(n3113), .B(n3737), .Y(n500) );
  OR2X2 U3071 ( .A(A[152]), .B(B[152]), .Y(n491) );
  AND2X2 U3072 ( .A(B[153]), .B(A[153]), .Y(n487) );
  INVX1 U3073 ( .A(n487), .Y(n3114) );
  OR2X1 U3074 ( .A(A[153]), .B(B[153]), .Y(n486) );
  INVX1 U3075 ( .A(n486), .Y(n3115) );
  OR2X2 U3076 ( .A(n502), .B(n482), .Y(n480) );
  INVX1 U3077 ( .A(n480), .Y(n3116) );
  OR2X2 U3078 ( .A(A[154]), .B(B[154]), .Y(n471) );
  OR2X1 U3079 ( .A(A[155]), .B(B[155]), .Y(n466) );
  OR2X2 U3080 ( .A(n4611), .B(n4516), .Y(n464) );
  INVX1 U3081 ( .A(n464), .Y(n3117) );
  AND2X2 U3082 ( .A(n584), .B(n4273), .Y(n454) );
  INVX1 U3083 ( .A(n454), .Y(n3118) );
  AND2X2 U3084 ( .A(B[156]), .B(A[156]), .Y(n450) );
  AND2X2 U3085 ( .A(B[157]), .B(A[157]), .Y(n443) );
  INVX1 U3086 ( .A(n443), .Y(n3119) );
  OR2X2 U3087 ( .A(n2953), .B(n3917), .Y(n438) );
  INVX1 U3088 ( .A(n438), .Y(n3120) );
  OR2X2 U3089 ( .A(n502), .B(n4312), .Y(n434) );
  INVX1 U3090 ( .A(n434), .Y(n3121) );
  OR2X2 U3091 ( .A(A[158]), .B(B[158]), .Y(n425) );
  AND2X2 U3092 ( .A(B[159]), .B(A[159]), .Y(n421) );
  INVX1 U3093 ( .A(n421), .Y(n3122) );
  OR2X1 U3094 ( .A(A[159]), .B(B[159]), .Y(n420) );
  AND2X2 U3095 ( .A(n4596), .B(n2945), .Y(n412) );
  INVX1 U3096 ( .A(n412), .Y(n3123) );
  OR2X2 U3097 ( .A(A[160]), .B(B[160]), .Y(n401) );
  OR2X2 U3098 ( .A(A[161]), .B(B[161]), .Y(n396) );
  OR2X2 U3099 ( .A(n4615), .B(n4521), .Y(n392) );
  INVX1 U3100 ( .A(n392), .Y(n3124) );
  OR2X2 U3101 ( .A(A[162]), .B(B[162]), .Y(n383) );
  OR2X2 U3102 ( .A(n3349), .B(n4618), .Y(n381) );
  INVX1 U3103 ( .A(n381), .Y(n3125) );
  AND2X2 U3104 ( .A(B[163]), .B(A[163]), .Y(n379) );
  INVX1 U3105 ( .A(n379), .Y(n3126) );
  OR2X2 U3106 ( .A(A[163]), .B(B[163]), .Y(n378) );
  OR2X2 U3107 ( .A(A[164]), .B(B[164]), .Y(n359) );
  INVX1 U3108 ( .A(n359), .Y(n3127) );
  OR2X2 U3109 ( .A(n3351), .B(n3127), .Y(n357) );
  INVX1 U3110 ( .A(n357), .Y(n3128) );
  AND2X2 U3111 ( .A(B[165]), .B(A[165]), .Y(n355) );
  INVX1 U3112 ( .A(n355), .Y(n3129) );
  OR2X2 U3113 ( .A(A[165]), .B(B[165]), .Y(n354) );
  OR2X2 U3114 ( .A(n4162), .B(n4619), .Y(n352) );
  OR2X2 U3115 ( .A(A[166]), .B(B[166]), .Y(n339) );
  OR2X2 U3116 ( .A(n3353), .B(n4622), .Y(n337) );
  INVX1 U3117 ( .A(n337), .Y(n3130) );
  AND2X2 U3118 ( .A(B[167]), .B(A[167]), .Y(n335) );
  INVX1 U3119 ( .A(n335), .Y(n3131) );
  OR2X2 U3120 ( .A(A[167]), .B(B[167]), .Y(n334) );
  INVX1 U3121 ( .A(n334), .Y(n3132) );
  OR2X2 U3122 ( .A(n3355), .B(n3463), .Y(n324) );
  OR2X2 U3123 ( .A(A[168]), .B(B[168]), .Y(n315) );
  OR2X2 U3124 ( .A(n3357), .B(n4624), .Y(n313) );
  INVX1 U3125 ( .A(n313), .Y(n3133) );
  AND2X2 U3126 ( .A(B[169]), .B(A[169]), .Y(n311) );
  INVX1 U3127 ( .A(n311), .Y(n3134) );
  OR2X2 U3128 ( .A(A[169]), .B(B[169]), .Y(n310) );
  AND2X2 U3129 ( .A(B[170]), .B(A[170]), .Y(n298) );
  OR2X2 U3130 ( .A(A[170]), .B(B[170]), .Y(n295) );
  OR2X2 U3131 ( .A(n3359), .B(n4625), .Y(n293) );
  INVX1 U3132 ( .A(n293), .Y(n3135) );
  AND2X2 U3133 ( .A(B[171]), .B(A[171]), .Y(n291) );
  INVX1 U3134 ( .A(n291), .Y(n3136) );
  OR2X2 U3135 ( .A(A[171]), .B(B[171]), .Y(n290) );
  AND2X2 U3136 ( .A(n3169), .B(n3563), .Y(n282) );
  OR2X2 U3137 ( .A(A[172]), .B(B[172]), .Y(n271) );
  OR2X2 U3138 ( .A(n3361), .B(n4630), .Y(n269) );
  INVX1 U3139 ( .A(n269), .Y(n3137) );
  OR2X2 U3140 ( .A(n4629), .B(n2954), .Y(n262) );
  INVX1 U3141 ( .A(n262), .Y(n3138) );
  AND2X2 U3142 ( .A(B[174]), .B(A[174]), .Y(n252) );
  OR2X2 U3143 ( .A(A[174]), .B(B[174]), .Y(n249) );
  OR2X2 U3144 ( .A(n3179), .B(n4631), .Y(n247) );
  INVX1 U3145 ( .A(n247), .Y(n3139) );
  AND2X2 U3146 ( .A(B[175]), .B(A[175]), .Y(n245) );
  INVX1 U3147 ( .A(n245), .Y(n3140) );
  OR2X2 U3148 ( .A(A[175]), .B(B[175]), .Y(n244) );
  OR2X2 U3149 ( .A(A[176]), .B(B[176]), .Y(n225) );
  INVX1 U3150 ( .A(n225), .Y(n3141) );
  OR2X2 U3151 ( .A(n3327), .B(n4633), .Y(n223) );
  INVX1 U3152 ( .A(n223), .Y(n3142) );
  AND2X2 U3153 ( .A(B[177]), .B(A[177]), .Y(n221) );
  INVX1 U3154 ( .A(n221), .Y(n3143) );
  OR2X2 U3155 ( .A(A[177]), .B(B[177]), .Y(n220) );
  OR2X2 U3156 ( .A(n3173), .B(n216), .Y(n214) );
  INVX1 U3157 ( .A(n214), .Y(n3144) );
  INVX1 U3158 ( .A(n352), .Y(n3145) );
  INVX1 U3159 ( .A(n484), .Y(n3146) );
  BUFX2 U3160 ( .A(n2067), .Y(n3147) );
  BUFX2 U3161 ( .A(n2000), .Y(n3148) );
  BUFX2 U3162 ( .A(n1931), .Y(n3149) );
  BUFX2 U3163 ( .A(n1843), .Y(n3150) );
  BUFX2 U3164 ( .A(n1839), .Y(n3151) );
  BUFX2 U3165 ( .A(n1770), .Y(n3152) );
  BUFX2 U3166 ( .A(n1688), .Y(n3153) );
  BUFX2 U3167 ( .A(n1492), .Y(n3154) );
  BUFX2 U3168 ( .A(n1423), .Y(n3155) );
  BUFX2 U3169 ( .A(n1255), .Y(n3156) );
  BUFX2 U3170 ( .A(n1165), .Y(n3157) );
  BUFX2 U3171 ( .A(n1161), .Y(n3158) );
  BUFX2 U3172 ( .A(n1071), .Y(n3159) );
  BUFX2 U3173 ( .A(n850), .Y(n3160) );
  BUFX2 U3174 ( .A(n833), .Y(n3161) );
  BUFX2 U3175 ( .A(n820), .Y(n3162) );
  BUFX2 U3176 ( .A(n803), .Y(n3163) );
  BUFX2 U3177 ( .A(n790), .Y(n3164) );
  BUFX2 U3178 ( .A(n773), .Y(n3165) );
  BUFX2 U3179 ( .A(n758), .Y(n3166) );
  BUFX2 U3180 ( .A(n741), .Y(n3167) );
  BUFX2 U3181 ( .A(n413), .Y(n3168) );
  OR2X2 U3182 ( .A(n4623), .B(n4526), .Y(n4138) );
  INVX1 U3183 ( .A(n4138), .Y(n3169) );
  INVX1 U3184 ( .A(n1676), .Y(n3170) );
  INVX1 U3185 ( .A(n1656), .Y(n3171) );
  INVX1 U3186 ( .A(n959), .Y(n3172) );
  INVX1 U3187 ( .A(n4321), .Y(n3173) );
  INVX1 U3188 ( .A(n4168), .Y(n3174) );
  INVX1 U3189 ( .A(n4747), .Y(n3175) );
  INVX1 U3190 ( .A(n4181), .Y(n3176) );
  INVX1 U3191 ( .A(n4702), .Y(n3177) );
  AND2X2 U3192 ( .A(n3117), .B(n3146), .Y(n458) );
  INVX1 U3193 ( .A(n458), .Y(n3178) );
  INVX1 U3194 ( .A(n4163), .Y(n3179) );
  OR2X2 U3195 ( .A(A[20]), .B(B[20]), .Y(n4144) );
  INVX1 U3196 ( .A(n4144), .Y(n3180) );
  AND2X2 U3197 ( .A(n3238), .B(n1966), .Y(n4145) );
  INVX1 U3198 ( .A(n4145), .Y(n3181) );
  OR2X2 U3199 ( .A(A[22]), .B(B[22]), .Y(n4146) );
  INVX1 U3200 ( .A(n4146), .Y(n3182) );
  INVX1 U3201 ( .A(n1791), .Y(n3183) );
  INVX1 U3202 ( .A(n1758), .Y(n3184) );
  INVX1 U3203 ( .A(n1740), .Y(n3185) );
  OR2X2 U3204 ( .A(A[46]), .B(B[46]), .Y(n4149) );
  INVX1 U3205 ( .A(n4149), .Y(n3186) );
  INVX1 U3206 ( .A(n1131), .Y(n3187) );
  INVX1 U3207 ( .A(n3752), .Y(n3188) );
  INVX1 U3208 ( .A(n827), .Y(n3189) );
  INVX1 U3209 ( .A(n4746), .Y(n3190) );
  INVX1 U3210 ( .A(n4692), .Y(n3191) );
  INVX1 U3211 ( .A(n4712), .Y(n3192) );
  OR2X2 U3212 ( .A(A[38]), .B(B[38]), .Y(n1780) );
  INVX1 U3213 ( .A(n4170), .Y(n3193) );
  INVX1 U3214 ( .A(n4762), .Y(n3194) );
  INVX1 U3215 ( .A(n4737), .Y(n3195) );
  INVX1 U3216 ( .A(n4715), .Y(n3196) );
  INVX1 U3217 ( .A(n4724), .Y(n3197) );
  INVX1 U3218 ( .A(n4771), .Y(n3198) );
  INVX1 U3219 ( .A(n4760), .Y(n3199) );
  OR2X2 U3220 ( .A(A[95]), .B(B[95]), .Y(n1168) );
  INVX1 U3221 ( .A(n1168), .Y(n3200) );
  INVX1 U3222 ( .A(n4736), .Y(n3201) );
  INVX1 U3223 ( .A(n4184), .Y(n3202) );
  OR2X2 U3224 ( .A(n3190), .B(n3604), .Y(n2095) );
  INVX1 U3225 ( .A(n2095), .Y(n3203) );
  INVX1 U3226 ( .A(n1179), .Y(n3204) );
  INVX1 U3227 ( .A(n4743), .Y(n3205) );
  INVX1 U3228 ( .A(n3741), .Y(n3206) );
  AND2X2 U3229 ( .A(n3315), .B(n3293), .Y(n2066) );
  INVX1 U3230 ( .A(n2066), .Y(n3207) );
  INVX1 U3231 ( .A(n3742), .Y(n3208) );
  AND2X2 U3232 ( .A(B[24]), .B(A[24]), .Y(n1922) );
  INVX1 U3233 ( .A(n1922), .Y(n3209) );
  AND2X2 U3234 ( .A(B[28]), .B(A[28]), .Y(n1880) );
  INVX1 U3235 ( .A(n1880), .Y(n3210) );
  INVX1 U3236 ( .A(n3745), .Y(n3211) );
  AND2X2 U3237 ( .A(B[60]), .B(A[60]), .Y(n1539) );
  INVX1 U3238 ( .A(n1539), .Y(n3212) );
  INVX1 U3239 ( .A(n3746), .Y(n3213) );
  INVX1 U3240 ( .A(n3747), .Y(n3214) );
  INVX1 U3241 ( .A(n3748), .Y(n3215) );
  AND2X2 U3242 ( .A(n2904), .B(n2895), .Y(n740) );
  INVX1 U3243 ( .A(n740), .Y(n3216) );
  AND2X2 U3244 ( .A(B[164]), .B(A[164]), .Y(n362) );
  INVX1 U3245 ( .A(n362), .Y(n3217) );
  INVX1 U3246 ( .A(n2114), .Y(n3218) );
  AND2X2 U3247 ( .A(B[72]), .B(A[72]), .Y(n4225) );
  INVX1 U3248 ( .A(n4225), .Y(n3219) );
  AND2X2 U3249 ( .A(B[96]), .B(A[96]), .Y(n4227) );
  INVX1 U3250 ( .A(n4227), .Y(n3220) );
  INVX1 U3251 ( .A(n4637), .Y(n3221) );
  INVX1 U3252 ( .A(n4754), .Y(n3222) );
  INVX1 U3253 ( .A(n3750), .Y(n3223) );
  INVX1 U3254 ( .A(n4692), .Y(n3224) );
  INVX1 U3255 ( .A(n4671), .Y(n3225) );
  INVX1 U3256 ( .A(n3743), .Y(n3226) );
  INVX1 U3257 ( .A(n4242), .Y(n3227) );
  AND2X2 U3258 ( .A(n4291), .B(n3295), .Y(n1838) );
  INVX1 U3259 ( .A(n1838), .Y(n3228) );
  INVX1 U3260 ( .A(n4480), .Y(n3229) );
  INVX1 U3261 ( .A(n4695), .Y(n3230) );
  BUFX2 U3262 ( .A(n237), .Y(n3231) );
  OR2X2 U3263 ( .A(A[67]), .B(B[67]), .Y(n4174) );
  INVX1 U3264 ( .A(n4174), .Y(n3232) );
  OR2X2 U3265 ( .A(A[100]), .B(B[100]), .Y(n4179) );
  INVX1 U3266 ( .A(n4179), .Y(n3233) );
  OR2X2 U3267 ( .A(A[124]), .B(B[124]), .Y(n4186) );
  INVX1 U3268 ( .A(n4186), .Y(n3234) );
  INVX1 U3269 ( .A(n4186), .Y(n3235) );
  OR2X2 U3270 ( .A(n3192), .B(n2873), .Y(n2001) );
  INVX1 U3271 ( .A(n2001), .Y(n3236) );
  OR2X2 U3272 ( .A(n3180), .B(n3410), .Y(n1948) );
  INVX1 U3273 ( .A(n1948), .Y(n3237) );
  INVX1 U3274 ( .A(n1948), .Y(n3238) );
  OR2X2 U3275 ( .A(n3887), .B(n3900), .Y(n1844) );
  INVX1 U3276 ( .A(n1844), .Y(n3239) );
  INVX1 U3277 ( .A(n1844), .Y(n3240) );
  OR2X2 U3278 ( .A(n3337), .B(n4481), .Y(n1551) );
  INVX1 U3279 ( .A(n1551), .Y(n3241) );
  OR2X2 U3280 ( .A(n3017), .B(n4453), .Y(n1497) );
  INVX1 U3281 ( .A(n1497), .Y(n3242) );
  INVX1 U3282 ( .A(n1497), .Y(n3243) );
  OR2X2 U3283 ( .A(n3342), .B(n3198), .Y(n1342) );
  INVX1 U3284 ( .A(n1342), .Y(n3244) );
  INVX1 U3285 ( .A(n1342), .Y(n3245) );
  OR2X2 U3286 ( .A(n3332), .B(n3408), .Y(n1982) );
  INVX1 U3287 ( .A(n1982), .Y(n3246) );
  OR2X2 U3288 ( .A(n3193), .B(n3407), .Y(n1707) );
  INVX1 U3289 ( .A(n1707), .Y(n3247) );
  INVX1 U3290 ( .A(n1707), .Y(n3248) );
  OR2X2 U3291 ( .A(n3232), .B(n3429), .Y(n1462) );
  INVX1 U3292 ( .A(n1462), .Y(n3249) );
  INVX1 U3293 ( .A(n1462), .Y(n3250) );
  OR2X2 U3294 ( .A(n3196), .B(n4488), .Y(n1276) );
  INVX1 U3295 ( .A(n1276), .Y(n3251) );
  INVX1 U3296 ( .A(n1276), .Y(n3252) );
  OR2X2 U3297 ( .A(n3189), .B(n4501), .Y(n812) );
  INVX1 U3298 ( .A(n812), .Y(n3253) );
  INVX1 U3299 ( .A(n812), .Y(n3254) );
  OR2X2 U3300 ( .A(n4372), .B(n4508), .Y(n552) );
  INVX1 U3301 ( .A(n552), .Y(n3255) );
  INVX1 U3302 ( .A(n552), .Y(n3256) );
  OR2X2 U3303 ( .A(n4613), .B(n4518), .Y(n418) );
  INVX1 U3304 ( .A(n418), .Y(n3257) );
  INVX1 U3305 ( .A(n418), .Y(n3258) );
  OR2X2 U3306 ( .A(n4620), .B(n3132), .Y(n332) );
  INVX1 U3307 ( .A(n332), .Y(n3259) );
  INVX1 U3308 ( .A(n332), .Y(n3260) );
  OR2X2 U3309 ( .A(n1866), .B(n4423), .Y(n1853) );
  INVX1 U3310 ( .A(n1853), .Y(n3261) );
  INVX1 U3311 ( .A(n1853), .Y(n3262) );
  OR2X2 U3312 ( .A(n3186), .B(n3421), .Y(n1689) );
  INVX1 U3313 ( .A(n1689), .Y(n3263) );
  INVX1 U3314 ( .A(n1689), .Y(n3264) );
  OR2X2 U3315 ( .A(n2855), .B(n4434), .Y(n1358) );
  INVX1 U3316 ( .A(n1358), .Y(n3265) );
  INVX1 U3317 ( .A(n1358), .Y(n3266) );
  OR2X2 U3318 ( .A(n670), .B(n4588), .Y(n624) );
  INVX1 U3319 ( .A(n624), .Y(n3267) );
  INVX1 U3320 ( .A(n624), .Y(n3268) );
  OR2X2 U3321 ( .A(n4167), .B(n3413), .Y(n2017) );
  INVX1 U3322 ( .A(n2017), .Y(n3269) );
  INVX1 U3323 ( .A(n2017), .Y(n3270) );
  OR2X2 U3324 ( .A(n3335), .B(n1787), .Y(n1785) );
  INVX1 U3325 ( .A(n1785), .Y(n3271) );
  INVX1 U3326 ( .A(n1785), .Y(n3272) );
  OR2X2 U3327 ( .A(n3184), .B(n3587), .Y(n1749) );
  INVX1 U3328 ( .A(n1749), .Y(n3273) );
  OR2X2 U3329 ( .A(n3733), .B(n3423), .Y(n1593) );
  INVX1 U3330 ( .A(n1593), .Y(n3274) );
  INVX1 U3331 ( .A(n1593), .Y(n3275) );
  OR2X2 U3332 ( .A(n3015), .B(n3425), .Y(n1521) );
  INVX1 U3333 ( .A(n1521), .Y(n3276) );
  INVX1 U3334 ( .A(n1521), .Y(n3277) );
  OR2X2 U3335 ( .A(n3341), .B(n3412), .Y(n1474) );
  INVX1 U3336 ( .A(n1474), .Y(n3278) );
  INVX1 U3337 ( .A(n1474), .Y(n3279) );
  OR2X2 U3338 ( .A(n3909), .B(n4153), .Y(n1232) );
  INVX1 U3339 ( .A(n1232), .Y(n3280) );
  INVX1 U3340 ( .A(n1232), .Y(n3281) );
  OR2X2 U3341 ( .A(n4600), .B(n4491), .Y(n1138) );
  INVX1 U3342 ( .A(n1138), .Y(n3282) );
  INVX1 U3343 ( .A(n1138), .Y(n3283) );
  OR2X2 U3344 ( .A(n3736), .B(n1092), .Y(n1090) );
  INVX1 U3345 ( .A(n1090), .Y(n3284) );
  OR2X2 U3346 ( .A(n4602), .B(n4499), .Y(n838) );
  INVX1 U3347 ( .A(n838), .Y(n3285) );
  INVX1 U3348 ( .A(n838), .Y(n3286) );
  OR2X2 U3349 ( .A(n4164), .B(n3141), .Y(n218) );
  INVX1 U3350 ( .A(n218), .Y(n3287) );
  AND2X2 U3351 ( .A(A[33]), .B(B[33]), .Y(n1832) );
  INVX1 U3352 ( .A(n1832), .Y(n3288) );
  OR2X2 U3353 ( .A(n3195), .B(n4486), .Y(n1316) );
  INVX1 U3354 ( .A(n1316), .Y(n3289) );
  INVX1 U3355 ( .A(n1316), .Y(n3290) );
  OR2X2 U3356 ( .A(n2914), .B(n3199), .Y(n1186) );
  INVX1 U3357 ( .A(n1186), .Y(n3291) );
  INVX1 U3358 ( .A(n1186), .Y(n3292) );
  OR2X2 U3359 ( .A(n3329), .B(n3411), .Y(n2080) );
  INVX1 U3360 ( .A(n2080), .Y(n3293) );
  INVX1 U3361 ( .A(n2080), .Y(n3294) );
  OR2X2 U3362 ( .A(n3498), .B(n3397), .Y(n1924) );
  INVX1 U3363 ( .A(n1924), .Y(n3295) );
  INVX1 U3364 ( .A(n1924), .Y(n3296) );
  OR2X2 U3365 ( .A(n3183), .B(n3418), .Y(n1789) );
  INVX1 U3366 ( .A(n1789), .Y(n3297) );
  INVX1 U3367 ( .A(n1789), .Y(n3298) );
  OR2X2 U3368 ( .A(n3194), .B(n4484), .Y(n1440) );
  INVX1 U3369 ( .A(n1440), .Y(n3299) );
  INVX1 U3370 ( .A(n1440), .Y(n3300) );
  OR2X2 U3371 ( .A(n4317), .B(n3593), .Y(n1248) );
  INVX1 U3372 ( .A(n1248), .Y(n3301) );
  INVX1 U3373 ( .A(n1248), .Y(n3302) );
  OR2X2 U3374 ( .A(n3188), .B(n4495), .Y(n1046) );
  INVX1 U3375 ( .A(n1046), .Y(n3303) );
  OR2X2 U3376 ( .A(n1064), .B(n4579), .Y(n1016) );
  INVX1 U3377 ( .A(n1016), .Y(n3304) );
  INVX1 U3378 ( .A(n1016), .Y(n3305) );
  OR2X2 U3379 ( .A(n1064), .B(n4306), .Y(n992) );
  INVX1 U3380 ( .A(n992), .Y(n3306) );
  OR2X2 U3381 ( .A(n4158), .B(n4505), .Y(n726) );
  INVX1 U3382 ( .A(n726), .Y(n3307) );
  INVX1 U3383 ( .A(n726), .Y(n3308) );
  OR2X2 U3384 ( .A(n4606), .B(n4510), .Y(n528) );
  INVX1 U3385 ( .A(n528), .Y(n3309) );
  INVX1 U3386 ( .A(n528), .Y(n3310) );
  OR2X2 U3387 ( .A(n3867), .B(n3200), .Y(n1166) );
  INVX1 U3388 ( .A(n1166), .Y(n3311) );
  INVX1 U3389 ( .A(n1166), .Y(n3312) );
  OR2X2 U3390 ( .A(n2883), .B(n3432), .Y(n1162) );
  INVX1 U3391 ( .A(n1162), .Y(n3313) );
  INVX1 U3392 ( .A(n1162), .Y(n3314) );
  OR2X2 U3393 ( .A(n3191), .B(n2877), .Y(n2068) );
  INVX1 U3394 ( .A(n2068), .Y(n3315) );
  INVX1 U3395 ( .A(n2068), .Y(n3316) );
  OR2X2 U3396 ( .A(n4157), .B(n4399), .Y(n924) );
  INVX1 U3397 ( .A(n924), .Y(n3317) );
  INVX1 U3398 ( .A(n924), .Y(n3318) );
  OR2X2 U3399 ( .A(n3197), .B(n3094), .Y(n714) );
  INVX1 U3400 ( .A(n714), .Y(n3319) );
  INVX1 U3401 ( .A(n714), .Y(n3320) );
  OR2X2 U3402 ( .A(n3905), .B(n4512), .Y(n508) );
  INVX1 U3403 ( .A(n508), .Y(n3321) );
  INVX1 U3404 ( .A(n508), .Y(n3322) );
  OR2X2 U3405 ( .A(n4609), .B(n3115), .Y(n484) );
  INVX1 U3406 ( .A(n484), .Y(n3323) );
  AND2X2 U3407 ( .A(n4279), .B(n4533), .Y(n1378) );
  INVX1 U3408 ( .A(n1378), .Y(n3324) );
  INVX1 U3409 ( .A(n1378), .Y(n3325) );
  AND2X2 U3410 ( .A(n3728), .B(n3052), .Y(n964) );
  INVX1 U3411 ( .A(n964), .Y(n3326) );
  AND2X2 U3412 ( .A(n234), .B(n406), .Y(n4321) );
  INVX1 U3413 ( .A(n4321), .Y(n3327) );
  INVX1 U3414 ( .A(n4321), .Y(n3328) );
  OR2X2 U3415 ( .A(A[4]), .B(B[4]), .Y(n2091) );
  INVX1 U3416 ( .A(n2091), .Y(n3329) );
  AND2X2 U3417 ( .A(n3730), .B(n2862), .Y(n2033) );
  INVX1 U3418 ( .A(n2033), .Y(n3330) );
  INVX1 U3419 ( .A(n2033), .Y(n3331) );
  OR2X2 U3420 ( .A(A[16]), .B(B[16]), .Y(n1993) );
  INVX1 U3421 ( .A(n1993), .Y(n3332) );
  AND2X2 U3422 ( .A(n2978), .B(n3721), .Y(n1884) );
  INVX1 U3423 ( .A(n1884), .Y(n3333) );
  INVX1 U3424 ( .A(n1884), .Y(n3334) );
  AND2X2 U3425 ( .A(n3567), .B(n4314), .Y(n1805) );
  INVX1 U3426 ( .A(n1805), .Y(n3335) );
  AND2X2 U3427 ( .A(n4532), .B(n1643), .Y(n1619) );
  INVX1 U3428 ( .A(n1619), .Y(n3336) );
  OR2X2 U3429 ( .A(A[58]), .B(B[58]), .Y(n1564) );
  INVX1 U3430 ( .A(n1564), .Y(n3337) );
  INVX1 U3431 ( .A(n1564), .Y(n3338) );
  AND2X2 U3432 ( .A(n3241), .B(n3723), .Y(n1545) );
  INVX1 U3433 ( .A(n1545), .Y(n3339) );
  INVX1 U3434 ( .A(n1545), .Y(n3340) );
  OR2X2 U3435 ( .A(A[64]), .B(B[64]), .Y(n1485) );
  INVX1 U3436 ( .A(n1485), .Y(n3341) );
  OR2X2 U3437 ( .A(A[79]), .B(B[79]), .Y(n1344) );
  INVX1 U3438 ( .A(n1344), .Y(n3342) );
  INVX1 U3439 ( .A(n1344), .Y(n3343) );
  OR2X2 U3440 ( .A(A[111]), .B(B[111]), .Y(n976) );
  INVX1 U3441 ( .A(n976), .Y(n3344) );
  INVX1 U3442 ( .A(n976), .Y(n3345) );
  AND2X2 U3443 ( .A(n4538), .B(n918), .Y(n892) );
  INVX1 U3444 ( .A(n892), .Y(n3346) );
  AND2X2 U3445 ( .A(n3253), .B(n3285), .Y(n806) );
  INVX1 U3446 ( .A(n806), .Y(n3347) );
  INVX1 U3447 ( .A(n806), .Y(n3348) );
  AND2X2 U3448 ( .A(n4547), .B(n406), .Y(n390) );
  INVX1 U3449 ( .A(n390), .Y(n3349) );
  INVX1 U3450 ( .A(n390), .Y(n3350) );
  AND2X2 U3451 ( .A(n368), .B(n406), .Y(n366) );
  INVX1 U3452 ( .A(n366), .Y(n3351) );
  INVX1 U3453 ( .A(n366), .Y(n3352) );
  AND2X2 U3454 ( .A(n2947), .B(n406), .Y(n346) );
  INVX1 U3455 ( .A(n346), .Y(n3353) );
  INVX1 U3456 ( .A(n346), .Y(n3354) );
  AND2X2 U3457 ( .A(n3259), .B(n3145), .Y(n330) );
  INVX1 U3458 ( .A(n330), .Y(n3355) );
  INVX1 U3459 ( .A(n330), .Y(n3356) );
  AND2X2 U3460 ( .A(n4599), .B(n406), .Y(n322) );
  INVX1 U3461 ( .A(n322), .Y(n3357) );
  INVX1 U3462 ( .A(n322), .Y(n3358) );
  AND2X2 U3463 ( .A(n2948), .B(n406), .Y(n302) );
  INVX1 U3464 ( .A(n302), .Y(n3359) );
  INVX1 U3465 ( .A(n302), .Y(n3360) );
  AND2X2 U3466 ( .A(n4287), .B(n406), .Y(n278) );
  INVX1 U3467 ( .A(n278), .Y(n3361) );
  INVX1 U3468 ( .A(n278), .Y(n3362) );
  AND2X2 U3469 ( .A(n3571), .B(n4598), .Y(n236) );
  INVX1 U3470 ( .A(n236), .Y(n3363) );
  INVX1 U3471 ( .A(n236), .Y(n3364) );
  AND2X2 U3472 ( .A(B[173]), .B(A[173]), .Y(n267) );
  INVX1 U3473 ( .A(n267), .Y(n3365) );
  AND2X2 U3474 ( .A(n4281), .B(n2848), .Y(n4152) );
  INVX1 U3475 ( .A(n4152), .Y(n3366) );
  INVX1 U3476 ( .A(n4152), .Y(n3367) );
  OR2X2 U3477 ( .A(A[10]), .B(B[10]), .Y(n2048) );
  OR2X2 U3478 ( .A(A[34]), .B(B[34]), .Y(n1820) );
  INVX1 U3479 ( .A(n1820), .Y(n3368) );
  INVX1 U3480 ( .A(n1820), .Y(n3369) );
  AND2X2 U3481 ( .A(n3247), .B(n3263), .Y(n1687) );
  INVX1 U3482 ( .A(n1687), .Y(n3370) );
  AND2X2 U3483 ( .A(n4534), .B(n2884), .Y(n1396) );
  INVX1 U3484 ( .A(n1396), .Y(n3371) );
  INVX1 U3485 ( .A(n1396), .Y(n3372) );
  AND2X2 U3486 ( .A(n3266), .B(n3025), .Y(n1356) );
  INVX1 U3487 ( .A(n1356), .Y(n3373) );
  INVX1 U3488 ( .A(n1356), .Y(n3374) );
  AND2X2 U3489 ( .A(n3290), .B(n2848), .Y(n1314) );
  INVX1 U3490 ( .A(n1314), .Y(n3375) );
  INVX1 U3491 ( .A(n1314), .Y(n3376) );
  AND2X2 U3492 ( .A(n4769), .B(n2848), .Y(n1246) );
  INVX1 U3493 ( .A(n1246), .Y(n3377) );
  INVX1 U3494 ( .A(n1246), .Y(n3378) );
  AND2X2 U3495 ( .A(n3068), .B(n3064), .Y(n972) );
  INVX1 U3496 ( .A(n972), .Y(n3379) );
  INVX1 U3497 ( .A(n972), .Y(n3380) );
  AND2X2 U3498 ( .A(n4540), .B(n708), .Y(n690) );
  INVX1 U3499 ( .A(n690), .Y(n3381) );
  INVX1 U3500 ( .A(n690), .Y(n3382) );
  AND2X2 U3501 ( .A(n4542), .B(n4590), .Y(n648) );
  INVX1 U3502 ( .A(n648), .Y(n3383) );
  INVX1 U3503 ( .A(n648), .Y(n3384) );
  AND2X2 U3504 ( .A(n4543), .B(n3267), .Y(n608) );
  INVX1 U3505 ( .A(n608), .Y(n3385) );
  INVX1 U3506 ( .A(n608), .Y(n3386) );
  AND2X2 U3507 ( .A(n4544), .B(n584), .Y(n566) );
  INVX1 U3508 ( .A(n566), .Y(n3387) );
  INVX1 U3509 ( .A(n566), .Y(n3388) );
  AND2X2 U3510 ( .A(n544), .B(n584), .Y(n542) );
  INVX1 U3511 ( .A(n542), .Y(n3389) );
  INVX1 U3512 ( .A(n542), .Y(n3390) );
  AND2X2 U3513 ( .A(n2943), .B(n584), .Y(n522) );
  INVX1 U3514 ( .A(n522), .Y(n3391) );
  INVX1 U3515 ( .A(n522), .Y(n3392) );
  AND2X2 U3516 ( .A(n4549), .B(n282), .Y(n260) );
  INVX1 U3517 ( .A(n260), .Y(n3393) );
  INVX1 U3518 ( .A(n260), .Y(n3394) );
  OR2X2 U3519 ( .A(A[56]), .B(B[56]), .Y(n1586) );
  INVX1 U3520 ( .A(n1586), .Y(n3395) );
  INVX1 U3521 ( .A(n1586), .Y(n3396) );
  AND2X2 U3522 ( .A(n3246), .B(n4700), .Y(n1964) );
  INVX1 U3523 ( .A(n1964), .Y(n3397) );
  INVX1 U3524 ( .A(n1964), .Y(n3398) );
  AND2X2 U3525 ( .A(n4141), .B(n2884), .Y(n1332) );
  INVX1 U3526 ( .A(n2848), .Y(n3399) );
  OR2X2 U3527 ( .A(A[83]), .B(B[83]), .Y(n1302) );
  INVX1 U3528 ( .A(n1302), .Y(n3400) );
  INVX1 U3529 ( .A(n1302), .Y(n3401) );
  AND2X2 U3530 ( .A(n4285), .B(n4594), .Y(n748) );
  INVX1 U3531 ( .A(n748), .Y(n3402) );
  INVX1 U3532 ( .A(n2907), .Y(n3403) );
  OR2X2 U3533 ( .A(A[27]), .B(B[27]), .Y(n4169) );
  INVX1 U3534 ( .A(n4169), .Y(n3404) );
  INVX1 U3535 ( .A(n4169), .Y(n3405) );
  OR2X2 U3536 ( .A(A[45]), .B(B[45]), .Y(n4171) );
  INVX1 U3537 ( .A(n4171), .Y(n3406) );
  INVX1 U3538 ( .A(n4171), .Y(n3407) );
  OR2X2 U3539 ( .A(A[17]), .B(B[17]), .Y(n4634) );
  INVX1 U3540 ( .A(n4634), .Y(n3408) );
  INVX1 U3541 ( .A(n4634), .Y(n3409) );
  OR2X2 U3542 ( .A(A[21]), .B(B[21]), .Y(n4637) );
  INVX1 U3543 ( .A(n4637), .Y(n3410) );
  OR2X2 U3544 ( .A(A[5]), .B(B[5]), .Y(n4671) );
  INVX1 U3545 ( .A(n4671), .Y(n3411) );
  OR2X2 U3546 ( .A(A[65]), .B(B[65]), .Y(n4695) );
  INVX1 U3547 ( .A(n4695), .Y(n3412) );
  OR2X2 U3548 ( .A(A[12]), .B(B[12]), .Y(n2030) );
  INVX1 U3549 ( .A(n2030), .Y(n3413) );
  INVX1 U3550 ( .A(n2030), .Y(n3414) );
  AND2X2 U3551 ( .A(n3239), .B(n2908), .Y(n1842) );
  INVX1 U3552 ( .A(n1842), .Y(n3415) );
  INVX1 U3553 ( .A(n1842), .Y(n3416) );
  OR2X2 U3554 ( .A(A[32]), .B(B[32]), .Y(n1834) );
  INVX1 U3555 ( .A(n1834), .Y(n3417) );
  OR2X2 U3556 ( .A(A[36]), .B(B[36]), .Y(n1798) );
  INVX1 U3557 ( .A(n1798), .Y(n3418) );
  INVX1 U3558 ( .A(n1798), .Y(n3419) );
  OR2X2 U3559 ( .A(A[39]), .B(B[39]), .Y(n1773) );
  INVX1 U3560 ( .A(n1773), .Y(n3420) );
  OR2X2 U3561 ( .A(A[47]), .B(B[47]), .Y(n1691) );
  INVX1 U3562 ( .A(n1691), .Y(n3421) );
  INVX1 U3563 ( .A(n1691), .Y(n3422) );
  AND2X2 U3564 ( .A(n2878), .B(n4531), .Y(n1599) );
  INVX1 U3565 ( .A(n1599), .Y(n3423) );
  INVX1 U3566 ( .A(n1599), .Y(n3424) );
  OR2X2 U3567 ( .A(A[60]), .B(B[60]), .Y(n1538) );
  INVX1 U3568 ( .A(n1538), .Y(n3425) );
  INVX1 U3569 ( .A(n1538), .Y(n3426) );
  AND2X2 U3570 ( .A(n3242), .B(n3276), .Y(n1495) );
  INVX1 U3571 ( .A(n1495), .Y(n3427) );
  INVX1 U3572 ( .A(n1495), .Y(n3428) );
  OR2X2 U3573 ( .A(A[66]), .B(B[66]), .Y(n1469) );
  INVX1 U3574 ( .A(n1469), .Y(n3429) );
  INVX1 U3575 ( .A(n1469), .Y(n3430) );
  AND2X2 U3576 ( .A(n2903), .B(n3280), .Y(n1206) );
  INVX1 U3577 ( .A(n1206), .Y(n3431) );
  INVX1 U3578 ( .A(n1206), .Y(n3432) );
  OR2X2 U3579 ( .A(A[103]), .B(B[103]), .Y(n1074) );
  INVX1 U3580 ( .A(n1074), .Y(n3433) );
  INVX1 U3581 ( .A(n1074), .Y(n3434) );
  OR2X2 U3582 ( .A(A[113]), .B(B[113]), .Y(n950) );
  INVX1 U3583 ( .A(n950), .Y(n3435) );
  INVX1 U3584 ( .A(n950), .Y(n3436) );
  AND2X2 U3585 ( .A(n2935), .B(n4689), .Y(n931) );
  INVX1 U3586 ( .A(n931), .Y(n3437) );
  INVX1 U3587 ( .A(n931), .Y(n3438) );
  AND2X2 U3588 ( .A(n918), .B(n2879), .Y(n914) );
  INVX1 U3589 ( .A(n914), .Y(n3439) );
  INVX1 U3590 ( .A(n914), .Y(n3440) );
  AND2X2 U3591 ( .A(n2938), .B(n4689), .Y(n903) );
  INVX1 U3592 ( .A(n903), .Y(n3441) );
  INVX1 U3593 ( .A(n903), .Y(n3442) );
  AND2X2 U3594 ( .A(n890), .B(n2879), .Y(n888) );
  INVX1 U3595 ( .A(n888), .Y(n3443) );
  AND2X2 U3596 ( .A(n3078), .B(n4689), .Y(n877) );
  INVX1 U3597 ( .A(n877), .Y(n3444) );
  INVX1 U3598 ( .A(n877), .Y(n3445) );
  AND2X2 U3599 ( .A(n4636), .B(n2879), .Y(n860) );
  INVX1 U3600 ( .A(n860), .Y(n3446) );
  INVX1 U3601 ( .A(n860), .Y(n3447) );
  AND2X2 U3602 ( .A(n2879), .B(n4259), .Y(n849) );
  INVX1 U3603 ( .A(n849), .Y(n3448) );
  INVX1 U3604 ( .A(n849), .Y(n3449) );
  AND2X2 U3605 ( .A(n4689), .B(n4261), .Y(n832) );
  INVX1 U3606 ( .A(n832), .Y(n3450) );
  INVX1 U3607 ( .A(n832), .Y(n3451) );
  AND2X2 U3608 ( .A(n2879), .B(n4263), .Y(n819) );
  INVX1 U3609 ( .A(n819), .Y(n3452) );
  INVX1 U3610 ( .A(n819), .Y(n3453) );
  AND2X2 U3611 ( .A(n4689), .B(n4265), .Y(n802) );
  INVX1 U3612 ( .A(n802), .Y(n3454) );
  INVX1 U3613 ( .A(n802), .Y(n3455) );
  AND2X2 U3614 ( .A(n4689), .B(n4267), .Y(n789) );
  INVX1 U3615 ( .A(n789), .Y(n3456) );
  INVX1 U3616 ( .A(n789), .Y(n3457) );
  AND2X2 U3617 ( .A(n4689), .B(n4269), .Y(n772) );
  INVX1 U3618 ( .A(n772), .Y(n3458) );
  INVX1 U3619 ( .A(n772), .Y(n3459) );
  AND2X2 U3620 ( .A(n2879), .B(n4271), .Y(n757) );
  INVX1 U3621 ( .A(n757), .Y(n3460) );
  INVX1 U3622 ( .A(n757), .Y(n3461) );
  AND2X2 U3623 ( .A(n3092), .B(n2846), .Y(n744) );
  INVX1 U3624 ( .A(n744), .Y(n3462) );
  AND2X2 U3625 ( .A(n3569), .B(n3124), .Y(n370) );
  INVX1 U3626 ( .A(n370), .Y(n3463) );
  INVX1 U3627 ( .A(n370), .Y(n3464) );
  BUFX2 U3628 ( .A(n1996), .Y(n3465) );
  AND2X2 U3629 ( .A(B[98]), .B(A[98]), .Y(n4213) );
  INVX1 U3630 ( .A(n4213), .Y(n3466) );
  INVX1 U3631 ( .A(n4213), .Y(n3467) );
  AND2X2 U3632 ( .A(B[50]), .B(A[50]), .Y(n4220) );
  INVX1 U3633 ( .A(n4220), .Y(n3468) );
  INVX1 U3634 ( .A(n4220), .Y(n3469) );
  AND2X2 U3635 ( .A(B[130]), .B(A[130]), .Y(n4228) );
  INVX1 U3636 ( .A(n4228), .Y(n3470) );
  INVX1 U3637 ( .A(n4228), .Y(n3471) );
  AND2X2 U3638 ( .A(B[64]), .B(A[64]), .Y(n1486) );
  INVX1 U3639 ( .A(n1486), .Y(n3472) );
  INVX1 U3640 ( .A(n1486), .Y(n3473) );
  AND2X2 U3641 ( .A(B[80]), .B(A[80]), .Y(n1328) );
  INVX1 U3642 ( .A(n1328), .Y(n3474) );
  INVX1 U3643 ( .A(n1328), .Y(n3475) );
  AND2X2 U3644 ( .A(B[88]), .B(A[88]), .Y(n1242) );
  INVX1 U3645 ( .A(n1242), .Y(n3476) );
  INVX1 U3646 ( .A(n1242), .Y(n3477) );
  AND2X2 U3647 ( .A(B[116]), .B(A[116]), .Y(n910) );
  INVX1 U3648 ( .A(n910), .Y(n3478) );
  INVX1 U3649 ( .A(n910), .Y(n3479) );
  AND2X2 U3650 ( .A(B[120]), .B(A[120]), .Y(n856) );
  INVX1 U3651 ( .A(n856), .Y(n3480) );
  INVX1 U3652 ( .A(n856), .Y(n3481) );
  AND2X2 U3653 ( .A(B[138]), .B(A[138]), .Y(n644) );
  INVX1 U3654 ( .A(n644), .Y(n3482) );
  INVX1 U3655 ( .A(n644), .Y(n3483) );
  AND2X2 U3656 ( .A(B[140]), .B(A[140]), .Y(n622) );
  INVX1 U3657 ( .A(n622), .Y(n3484) );
  INVX1 U3658 ( .A(n622), .Y(n3485) );
  AND2X2 U3659 ( .A(B[142]), .B(A[142]), .Y(n604) );
  INVX1 U3660 ( .A(n604), .Y(n3486) );
  INVX1 U3661 ( .A(n604), .Y(n3487) );
  AND2X2 U3662 ( .A(B[162]), .B(A[162]), .Y(n386) );
  INVX1 U3663 ( .A(n386), .Y(n3488) );
  INVX1 U3664 ( .A(n386), .Y(n3489) );
  AND2X2 U3665 ( .A(B[168]), .B(A[168]), .Y(n318) );
  INVX1 U3666 ( .A(n318), .Y(n3490) );
  INVX1 U3667 ( .A(n318), .Y(n3491) );
  AND2X2 U3668 ( .A(B[176]), .B(A[176]), .Y(n228) );
  INVX1 U3669 ( .A(n228), .Y(n3492) );
  INVX1 U3670 ( .A(n228), .Y(n3493) );
  AND2X2 U3671 ( .A(B[2]), .B(A[2]), .Y(n2101) );
  INVX1 U3672 ( .A(n2101), .Y(n3494) );
  INVX1 U3673 ( .A(n2101), .Y(n3495) );
  AND2X2 U3674 ( .A(B[8]), .B(A[8]), .Y(n2063) );
  INVX1 U3675 ( .A(n2063), .Y(n3496) );
  INVX1 U3676 ( .A(n2063), .Y(n3497) );
  AND2X2 U3677 ( .A(n3237), .B(n3565), .Y(n1930) );
  INVX1 U3678 ( .A(n1930), .Y(n3498) );
  AND2X2 U3679 ( .A(B[42]), .B(A[42]), .Y(n1741) );
  INVX1 U3680 ( .A(n1741), .Y(n3499) );
  BUFX2 U3681 ( .A(n2094), .Y(n3500) );
  BUFX2 U3682 ( .A(n2034), .Y(n3501) );
  BUFX2 U3683 ( .A(n1806), .Y(n3502) );
  BUFX2 U3684 ( .A(n1457), .Y(n3503) );
  BUFX2 U3685 ( .A(n1381), .Y(n3504) );
  BUFX2 U3686 ( .A(n1333), .Y(n3505) );
  BUFX2 U3687 ( .A(n633), .Y(n3506) );
  AND2X2 U3688 ( .A(B[70]), .B(A[70]), .Y(n4224) );
  INVX1 U3689 ( .A(n4224), .Y(n3507) );
  INVX1 U3690 ( .A(n4224), .Y(n3508) );
  AND2X2 U3691 ( .A(B[10]), .B(A[10]), .Y(n2049) );
  INVX1 U3692 ( .A(n2049), .Y(n3509) );
  INVX1 U3693 ( .A(n2049), .Y(n3510) );
  AND2X2 U3694 ( .A(B[14]), .B(A[14]), .Y(n2013) );
  INVX1 U3695 ( .A(n2013), .Y(n3511) );
  INVX1 U3696 ( .A(n2013), .Y(n3512) );
  AND2X2 U3697 ( .A(B[32]), .B(A[32]), .Y(n1835) );
  INVX1 U3698 ( .A(n1835), .Y(n3513) );
  INVX1 U3699 ( .A(n1835), .Y(n3514) );
  AND2X2 U3700 ( .A(B[76]), .B(A[76]), .Y(n1370) );
  INVX1 U3701 ( .A(n1370), .Y(n3515) );
  INVX1 U3702 ( .A(n1370), .Y(n3516) );
  AND2X2 U3703 ( .A(B[118]), .B(A[118]), .Y(n884) );
  INVX1 U3704 ( .A(n884), .Y(n3517) );
  INVX1 U3705 ( .A(n884), .Y(n3518) );
  AND2X2 U3706 ( .A(B[126]), .B(A[126]), .Y(n768) );
  INVX1 U3707 ( .A(n768), .Y(n3519) );
  INVX1 U3708 ( .A(n768), .Y(n3520) );
  AND2X2 U3709 ( .A(B[136]), .B(A[136]), .Y(n662) );
  INVX1 U3710 ( .A(n662), .Y(n3521) );
  INVX1 U3711 ( .A(n662), .Y(n3522) );
  AND2X2 U3712 ( .A(B[172]), .B(A[172]), .Y(n274) );
  INVX1 U3713 ( .A(n274), .Y(n3523) );
  INVX1 U3714 ( .A(n274), .Y(n3524) );
  BUFX2 U3715 ( .A(n1965), .Y(n3525) );
  BUFX2 U3716 ( .A(n1726), .Y(n3526) );
  BUFX2 U3717 ( .A(n1680), .Y(n3527) );
  BUFX2 U3718 ( .A(n1642), .Y(n3528) );
  BUFX2 U3719 ( .A(n1546), .Y(n3529) );
  BUFX2 U3720 ( .A(n1397), .Y(n3530) );
  BUFX2 U3721 ( .A(n1357), .Y(n3531) );
  BUFX2 U3722 ( .A(n1295), .Y(n3532) );
  BUFX2 U3723 ( .A(n1207), .Y(n3533) );
  BUFX2 U3724 ( .A(n1115), .Y(n3534) );
  BUFX2 U3725 ( .A(n1019), .Y(n3535) );
  BUFX2 U3726 ( .A(n919), .Y(n3536) );
  BUFX2 U3727 ( .A(n709), .Y(n3537) );
  BUFX2 U3728 ( .A(n649), .Y(n3538) );
  BUFX2 U3729 ( .A(n609), .Y(n3539) );
  BUFX2 U3730 ( .A(n585), .Y(n3540) );
  BUFX2 U3731 ( .A(n547), .Y(n3541) );
  BUFX2 U3732 ( .A(n479), .Y(n3542) );
  BUFX2 U3733 ( .A(n459), .Y(n3543) );
  BUFX2 U3734 ( .A(n455), .Y(n3544) );
  BUFX2 U3735 ( .A(n433), .Y(n3545) );
  BUFX2 U3736 ( .A(n391), .Y(n3546) );
  BUFX2 U3737 ( .A(n371), .Y(n3547) );
  BUFX2 U3738 ( .A(n367), .Y(n3548) );
  BUFX2 U3739 ( .A(n347), .Y(n3549) );
  BUFX2 U3740 ( .A(n323), .Y(n3550) );
  BUFX2 U3741 ( .A(n303), .Y(n3551) );
  BUFX2 U3742 ( .A(n279), .Y(n3552) );
  BUFX2 U3743 ( .A(n257), .Y(n3553) );
  BUFX2 U3744 ( .A(n233), .Y(n3554) );
  AND2X2 U3745 ( .A(B[34]), .B(A[34]), .Y(n1821) );
  INVX1 U3746 ( .A(n1821), .Y(n3555) );
  INVX1 U3747 ( .A(n1821), .Y(n3556) );
  OR2X2 U3748 ( .A(n3185), .B(n2996), .Y(n1731) );
  INVX1 U3749 ( .A(n1731), .Y(n3557) );
  INVX1 U3750 ( .A(n1731), .Y(n3558) );
  OR2X2 U3751 ( .A(n3187), .B(n3046), .Y(n1120) );
  INVX1 U3752 ( .A(n1120), .Y(n3559) );
  INVX1 U3753 ( .A(n1120), .Y(n3560) );
  OR2X2 U3754 ( .A(n4189), .B(n4631), .Y(n242) );
  INVX1 U3755 ( .A(n242), .Y(n3561) );
  INVX1 U3756 ( .A(n242), .Y(n3562) );
  OR2X2 U3757 ( .A(n4188), .B(n4625), .Y(n288) );
  INVX1 U3758 ( .A(n288), .Y(n3563) );
  INVX1 U3759 ( .A(n288), .Y(n3564) );
  OR2X2 U3760 ( .A(n3182), .B(n2971), .Y(n1932) );
  INVX1 U3761 ( .A(n1932), .Y(n3565) );
  INVX1 U3762 ( .A(n1932), .Y(n3566) );
  OR2X2 U3763 ( .A(n3368), .B(n3591), .Y(n1811) );
  INVX1 U3764 ( .A(n1811), .Y(n3567) );
  INVX1 U3765 ( .A(n1811), .Y(n3568) );
  OR2X2 U3766 ( .A(n4522), .B(n4617), .Y(n376) );
  INVX1 U3767 ( .A(n376), .Y(n3569) );
  INVX1 U3768 ( .A(n376), .Y(n3570) );
  OR2X2 U3769 ( .A(n4627), .B(n3601), .Y(n238) );
  INVX1 U3770 ( .A(n238), .Y(n3571) );
  INVX1 U3771 ( .A(n238), .Y(n3572) );
  AND2X2 U3772 ( .A(n4140), .B(n3274), .Y(n1491) );
  INVX1 U3773 ( .A(n1491), .Y(n3573) );
  INVX1 U3774 ( .A(n1491), .Y(n3574) );
  BUFX2 U3775 ( .A(n2088), .Y(n3575) );
  BUFX2 U3776 ( .A(n1943), .Y(n3576) );
  BUFX2 U3777 ( .A(n1903), .Y(n3577) );
  BUFX2 U3778 ( .A(n1894), .Y(n3578) );
  BUFX2 U3779 ( .A(n1133), .Y(n3579) );
  BUFX2 U3780 ( .A(n605), .Y(n3580) );
  BUFX2 U3781 ( .A(n539), .Y(n3581) );
  BUFX2 U3782 ( .A(n519), .Y(n3582) );
  BUFX2 U3783 ( .A(n468), .Y(n3583) );
  BUFX2 U3784 ( .A(n380), .Y(n3584) );
  BUFX2 U3785 ( .A(n343), .Y(n3585) );
  BUFX2 U3786 ( .A(n319), .Y(n3586) );
  OR2X2 U3787 ( .A(A[41]), .B(B[41]), .Y(n4477) );
  INVX1 U3788 ( .A(n4477), .Y(n3587) );
  OR2X2 U3789 ( .A(A[11]), .B(B[11]), .Y(n2041) );
  INVX1 U3790 ( .A(n2041), .Y(n3588) );
  AND2X2 U3791 ( .A(n3236), .B(n3269), .Y(n1999) );
  INVX1 U3792 ( .A(n1999), .Y(n3589) );
  INVX1 U3793 ( .A(n1999), .Y(n3590) );
  OR2X2 U3794 ( .A(A[35]), .B(B[35]), .Y(n1813) );
  INVX1 U3795 ( .A(n1813), .Y(n3591) );
  INVX1 U3796 ( .A(n1813), .Y(n3592) );
  AND2X2 U3797 ( .A(n3251), .B(n2886), .Y(n1254) );
  INVX1 U3798 ( .A(n1254), .Y(n3593) );
  INVX1 U3799 ( .A(n1254), .Y(n3594) );
  AND2X2 U3800 ( .A(n3051), .B(n2840), .Y(n1070) );
  INVX1 U3801 ( .A(n1070), .Y(n3595) );
  INVX1 U3802 ( .A(n1070), .Y(n3596) );
  AND2X2 U3803 ( .A(n3098), .B(n4539), .Y(n674) );
  INVX1 U3804 ( .A(n674), .Y(n3597) );
  INVX1 U3805 ( .A(n674), .Y(n3598) );
  AND2X2 U3806 ( .A(n3257), .B(n3120), .Y(n416) );
  INVX1 U3807 ( .A(n416), .Y(n3599) );
  INVX1 U3808 ( .A(n416), .Y(n3600) );
  AND2X2 U3809 ( .A(n3562), .B(n3138), .Y(n240) );
  INVX1 U3810 ( .A(n240), .Y(n3601) );
  INVX1 U3811 ( .A(n240), .Y(n3602) );
  OR2X2 U3812 ( .A(A[3]), .B(B[3]), .Y(n2097) );
  INVX1 U3813 ( .A(n2097), .Y(n3603) );
  INVX1 U3814 ( .A(n2097), .Y(n3604) );
  BUFX2 U3815 ( .A(n2079), .Y(n3605) );
  BUFX2 U3816 ( .A(n1990), .Y(n3606) );
  BUFX2 U3817 ( .A(n1961), .Y(n3607) );
  BUFX2 U3818 ( .A(n1954), .Y(n3608) );
  BUFX2 U3819 ( .A(n1936), .Y(n3609) );
  BUFX2 U3820 ( .A(n1923), .Y(n3610) );
  BUFX2 U3821 ( .A(n1916), .Y(n3611) );
  BUFX2 U3822 ( .A(n1881), .Y(n3612) );
  BUFX2 U3823 ( .A(n1872), .Y(n3613) );
  BUFX2 U3824 ( .A(n1859), .Y(n3614) );
  BUFX2 U3825 ( .A(n1482), .Y(n3615) );
  BUFX2 U3826 ( .A(n1473), .Y(n3616) );
  BUFX2 U3827 ( .A(n1466), .Y(n3617) );
  BUFX2 U3828 ( .A(n1453), .Y(n3618) );
  BUFX2 U3829 ( .A(n1446), .Y(n3619) );
  BUFX2 U3830 ( .A(n1435), .Y(n3620) );
  BUFX2 U3831 ( .A(n1428), .Y(n3621) );
  BUFX2 U3832 ( .A(n1411), .Y(n3622) );
  BUFX2 U3833 ( .A(n1404), .Y(n3623) );
  BUFX2 U3834 ( .A(n1393), .Y(n3624) );
  BUFX2 U3835 ( .A(n1386), .Y(n3625) );
  BUFX2 U3836 ( .A(n1371), .Y(n3626) );
  BUFX2 U3837 ( .A(n1364), .Y(n3627) );
  BUFX2 U3838 ( .A(n1353), .Y(n3628) );
  BUFX2 U3839 ( .A(n1346), .Y(n3629) );
  BUFX2 U3840 ( .A(n1329), .Y(n3630) );
  BUFX2 U3841 ( .A(n1322), .Y(n3631) );
  BUFX2 U3842 ( .A(n1311), .Y(n3632) );
  BUFX2 U3843 ( .A(n1304), .Y(n3633) );
  BUFX2 U3844 ( .A(n1287), .Y(n3634) );
  BUFX2 U3845 ( .A(n1280), .Y(n3635) );
  BUFX2 U3846 ( .A(n1267), .Y(n3636) );
  BUFX2 U3847 ( .A(n1260), .Y(n3637) );
  BUFX2 U3848 ( .A(n1243), .Y(n3638) );
  BUFX2 U3849 ( .A(n1236), .Y(n3639) );
  BUFX2 U3850 ( .A(n1223), .Y(n3640) );
  BUFX2 U3851 ( .A(n1216), .Y(n3641) );
  BUFX2 U3852 ( .A(n1199), .Y(n3642) );
  BUFX2 U3853 ( .A(n1192), .Y(n3643) );
  BUFX2 U3854 ( .A(n1177), .Y(n3644) );
  BUFX2 U3855 ( .A(n1170), .Y(n3645) );
  BUFX2 U3856 ( .A(n1153), .Y(n3646) );
  BUFX2 U3857 ( .A(n1146), .Y(n3647) );
  BUFX2 U3858 ( .A(n1124), .Y(n3648) );
  BUFX2 U3859 ( .A(n1107), .Y(n3649) );
  BUFX2 U3860 ( .A(n1098), .Y(n3650) );
  BUFX2 U3861 ( .A(n1085), .Y(n3651) );
  BUFX2 U3862 ( .A(n1076), .Y(n3652) );
  BUFX2 U3863 ( .A(n1059), .Y(n3653) );
  BUFX2 U3864 ( .A(n1050), .Y(n3654) );
  BUFX2 U3865 ( .A(n1037), .Y(n3655) );
  BUFX2 U3866 ( .A(n1028), .Y(n3656) );
  BUFX2 U3867 ( .A(n1011), .Y(n3657) );
  BUFX2 U3868 ( .A(n1002), .Y(n3658) );
  BUFX2 U3869 ( .A(n987), .Y(n3659) );
  BUFX2 U3870 ( .A(n978), .Y(n3660) );
  BUFX2 U3871 ( .A(n961), .Y(n3661) );
  BUFX2 U3872 ( .A(n952), .Y(n3662) );
  BUFX2 U3873 ( .A(n939), .Y(n3663) );
  BUFX2 U3874 ( .A(n928), .Y(n3664) );
  BUFX2 U3875 ( .A(n911), .Y(n3665) );
  BUFX2 U3876 ( .A(n900), .Y(n3666) );
  BUFX2 U3877 ( .A(n885), .Y(n3667) );
  BUFX2 U3878 ( .A(n874), .Y(n3668) );
  BUFX2 U3879 ( .A(n857), .Y(n3669) );
  BUFX2 U3880 ( .A(n846), .Y(n3670) );
  BUFX2 U3881 ( .A(n829), .Y(n3671) );
  BUFX2 U3882 ( .A(n816), .Y(n3672) );
  BUFX2 U3883 ( .A(n799), .Y(n3673) );
  BUFX2 U3884 ( .A(n786), .Y(n3674) );
  BUFX2 U3885 ( .A(n769), .Y(n3675) );
  BUFX2 U3886 ( .A(n754), .Y(n3676) );
  BUFX2 U3887 ( .A(n734), .Y(n3677) );
  BUFX2 U3888 ( .A(n725), .Y(n3678) );
  BUFX2 U3889 ( .A(n718), .Y(n3679) );
  BUFX2 U3890 ( .A(n705), .Y(n3680) );
  BUFX2 U3891 ( .A(n698), .Y(n3681) );
  BUFX2 U3892 ( .A(n687), .Y(n3682) );
  BUFX2 U3893 ( .A(n680), .Y(n3683) );
  BUFX2 U3894 ( .A(n663), .Y(n3684) );
  BUFX2 U3895 ( .A(n656), .Y(n3685) );
  BUFX2 U3896 ( .A(n645), .Y(n3686) );
  BUFX2 U3897 ( .A(n638), .Y(n3687) );
  BUFX2 U3898 ( .A(n623), .Y(n3688) );
  BUFX2 U3899 ( .A(n616), .Y(n3689) );
  BUFX2 U3900 ( .A(n598), .Y(n3690) );
  BUFX2 U3901 ( .A(n581), .Y(n3691) );
  BUFX2 U3902 ( .A(n574), .Y(n3692) );
  BUFX2 U3903 ( .A(n563), .Y(n3693) );
  BUFX2 U3904 ( .A(n556), .Y(n3694) );
  BUFX2 U3905 ( .A(n532), .Y(n3695) );
  BUFX2 U3906 ( .A(n512), .Y(n3696) );
  BUFX2 U3907 ( .A(n495), .Y(n3697) );
  BUFX2 U3908 ( .A(n488), .Y(n3698) );
  BUFX2 U3909 ( .A(n475), .Y(n3699) );
  BUFX2 U3910 ( .A(n451), .Y(n3700) );
  BUFX2 U3911 ( .A(n444), .Y(n3701) );
  BUFX2 U3912 ( .A(n429), .Y(n3702) );
  BUFX2 U3913 ( .A(n422), .Y(n3703) );
  BUFX2 U3914 ( .A(n405), .Y(n3704) );
  BUFX2 U3915 ( .A(n398), .Y(n3705) );
  BUFX2 U3916 ( .A(n387), .Y(n3706) );
  BUFX2 U3917 ( .A(n363), .Y(n3707) );
  BUFX2 U3918 ( .A(n356), .Y(n3708) );
  BUFX2 U3919 ( .A(n336), .Y(n3709) );
  BUFX2 U3920 ( .A(n312), .Y(n3710) );
  BUFX2 U3921 ( .A(n299), .Y(n3711) );
  BUFX2 U3922 ( .A(n292), .Y(n3712) );
  BUFX2 U3923 ( .A(n275), .Y(n3713) );
  BUFX2 U3924 ( .A(n268), .Y(n3714) );
  BUFX2 U3925 ( .A(n253), .Y(n3715) );
  BUFX2 U3926 ( .A(n246), .Y(n3716) );
  BUFX2 U3927 ( .A(n229), .Y(n3717) );
  BUFX2 U3928 ( .A(n222), .Y(n3718) );
  BUFX2 U3929 ( .A(n213), .Y(n3719) );
  BUFX2 U3930 ( .A(n200), .Y(n3720) );
  OR2X2 U3931 ( .A(n4147), .B(n3227), .Y(n1908) );
  INVX1 U3932 ( .A(n1908), .Y(n3721) );
  INVX1 U3933 ( .A(n1908), .Y(n3722) );
  OR2X2 U3934 ( .A(n4452), .B(n3395), .Y(n1573) );
  INVX1 U3935 ( .A(n1573), .Y(n3723) );
  INVX1 U3936 ( .A(n1573), .Y(n3724) );
  AND2X2 U3937 ( .A(n3558), .B(n3273), .Y(n1725) );
  INVX1 U3938 ( .A(n1725), .Y(n3725) );
  AND2X2 U3939 ( .A(n2912), .B(n2906), .Y(n1679) );
  INVX1 U3940 ( .A(n1679), .Y(n3726) );
  INVX1 U3941 ( .A(n1679), .Y(n3727) );
  OR2X2 U3942 ( .A(n3379), .B(n4578), .Y(n970) );
  INVX1 U3943 ( .A(n970), .Y(n3728) );
  INVX1 U3944 ( .A(n970), .Y(n3729) );
  OR2X2 U3945 ( .A(n2961), .B(n4679), .Y(n2053) );
  INVX1 U3946 ( .A(n2053), .Y(n3730) );
  INVX1 U3947 ( .A(n2053), .Y(n3731) );
  AND2X2 U3948 ( .A(n3495), .B(n4746), .Y(n195) );
  INVX1 U3949 ( .A(n195), .Y(n3732) );
  AND2X2 U3950 ( .A(n4139), .B(n4591), .Y(n1641) );
  INVX1 U3951 ( .A(n1641), .Y(n3733) );
  INVX1 U3952 ( .A(n1641), .Y(n3734) );
  AND2X2 U3953 ( .A(n3560), .B(n3282), .Y(n1114) );
  INVX1 U3954 ( .A(n1114), .Y(n3735) );
  INVX1 U3955 ( .A(n1114), .Y(n3736) );
  AND2X2 U3956 ( .A(n3255), .B(n3111), .Y(n546) );
  INVX1 U3957 ( .A(n546), .Y(n3737) );
  INVX1 U3958 ( .A(n546), .Y(n3738) );
  BUFX2 U3959 ( .A(n965), .Y(n3739) );
  AND2X2 U3960 ( .A(B[4]), .B(A[4]), .Y(n3741) );
  AND2X2 U3961 ( .A(B[12]), .B(A[12]), .Y(n3742) );
  AND2X2 U3962 ( .A(B[16]), .B(A[16]), .Y(n3743) );
  AND2X2 U3963 ( .A(B[48]), .B(A[48]), .Y(n3744) );
  AND2X2 U3964 ( .A(B[58]), .B(A[58]), .Y(n3745) );
  AND2X2 U3965 ( .A(B[104]), .B(A[104]), .Y(n3746) );
  AND2X2 U3966 ( .A(B[112]), .B(A[112]), .Y(n3747) );
  AND2X2 U3967 ( .A(B[124]), .B(A[124]), .Y(n3748) );
  OR2X2 U3968 ( .A(n2019), .B(n4403), .Y(n3749) );
  AND2X2 U3969 ( .A(B[40]), .B(A[40]), .Y(n3750) );
  AND2X2 U3970 ( .A(B[86]), .B(A[86]), .Y(n3751) );
  OR2X2 U3971 ( .A(A[104]), .B(B[104]), .Y(n3752) );
  OR2X2 U3972 ( .A(n4623), .B(n4527), .Y(n3753) );
  INVX1 U3973 ( .A(n4761), .Y(n3754) );
  BUFX2 U3974 ( .A(n2045), .Y(n3755) );
  INVX1 U3975 ( .A(n2027), .Y(n3756) );
  INVX1 U3976 ( .A(n3756), .Y(n3757) );
  INVX1 U3977 ( .A(n2016), .Y(n3758) );
  INVX1 U3978 ( .A(n3758), .Y(n3759) );
  INVX1 U3979 ( .A(n2007), .Y(n3760) );
  INVX1 U3980 ( .A(n3760), .Y(n3761) );
  BUFX2 U3981 ( .A(n1898), .Y(n3762) );
  BUFX2 U3982 ( .A(n1876), .Y(n3763) );
  BUFX2 U3983 ( .A(n1863), .Y(n3764) );
  BUFX2 U3984 ( .A(n1852), .Y(n3765) );
  BUFX2 U3985 ( .A(n1817), .Y(n3766) );
  BUFX2 U3986 ( .A(n1795), .Y(n3767) );
  BUFX2 U3987 ( .A(n1777), .Y(n3768) );
  BUFX2 U3988 ( .A(n1755), .Y(n3769) );
  BUFX2 U3989 ( .A(n1737), .Y(n3770) );
  BUFX2 U3990 ( .A(n1715), .Y(n3771) );
  BUFX2 U3991 ( .A(n1706), .Y(n3772) );
  BUFX2 U3992 ( .A(n1695), .Y(n3773) );
  INVX1 U3993 ( .A(n1673), .Y(n3774) );
  INVX1 U3994 ( .A(n3774), .Y(n3775) );
  INVX1 U3995 ( .A(n1662), .Y(n3776) );
  INVX1 U3996 ( .A(n3776), .Y(n3777) );
  INVX1 U3997 ( .A(n1653), .Y(n3778) );
  INVX1 U3998 ( .A(n3778), .Y(n3779) );
  INVX1 U3999 ( .A(n1638), .Y(n3780) );
  INVX1 U4000 ( .A(n3780), .Y(n3781) );
  INVX1 U4001 ( .A(n1629), .Y(n3782) );
  INVX1 U4002 ( .A(n3782), .Y(n3783) );
  INVX1 U4003 ( .A(n1616), .Y(n3784) );
  INVX1 U4004 ( .A(n3784), .Y(n3785) );
  INVX1 U4005 ( .A(n1607), .Y(n3786) );
  INVX1 U4006 ( .A(n3786), .Y(n3787) );
  INVX1 U4007 ( .A(n1600), .Y(n3788) );
  INVX1 U4008 ( .A(n3788), .Y(n3789) );
  INVX1 U4009 ( .A(n1592), .Y(n3790) );
  INVX1 U4010 ( .A(n3790), .Y(n3791) );
  INVX1 U4011 ( .A(n1583), .Y(n3792) );
  INVX1 U4012 ( .A(n3792), .Y(n3793) );
  INVX1 U4013 ( .A(n1568), .Y(n3794) );
  INVX1 U4014 ( .A(n3794), .Y(n3795) );
  BUFX2 U4015 ( .A(n1561), .Y(n3796) );
  INVX1 U4016 ( .A(n1557), .Y(n3797) );
  INVX1 U4017 ( .A(n3797), .Y(n3798) );
  INVX1 U4018 ( .A(n1542), .Y(n3799) );
  INVX1 U4019 ( .A(n3799), .Y(n3800) );
  BUFX2 U4020 ( .A(n1535), .Y(n3801) );
  INVX1 U4021 ( .A(n1531), .Y(n3802) );
  INVX1 U4022 ( .A(n3802), .Y(n3803) );
  BUFX2 U4023 ( .A(n1520), .Y(n3804) );
  INVX1 U4024 ( .A(n1516), .Y(n3805) );
  INVX1 U4025 ( .A(n3805), .Y(n3806) );
  BUFX2 U4026 ( .A(n1507), .Y(n3807) );
  INVX1 U4027 ( .A(n1503), .Y(n3808) );
  INVX1 U4028 ( .A(n3808), .Y(n3809) );
  INVX1 U4029 ( .A(n1496), .Y(n3810) );
  INVX1 U4030 ( .A(n3810), .Y(n3811) );
  INVX1 U4031 ( .A(n1341), .Y(n3812) );
  INVX1 U4032 ( .A(n3812), .Y(n3813) );
  INVX1 U4033 ( .A(n1185), .Y(n3814) );
  INVX1 U4034 ( .A(n3814), .Y(n3815) );
  BUFX2 U4035 ( .A(n1128), .Y(n3816) );
  BUFX2 U4036 ( .A(n1102), .Y(n3817) );
  BUFX2 U4037 ( .A(n1080), .Y(n3818) );
  BUFX2 U4038 ( .A(n1054), .Y(n3819) );
  BUFX2 U4039 ( .A(n1032), .Y(n3820) );
  INVX1 U4040 ( .A(n1006), .Y(n3821) );
  INVX1 U4041 ( .A(n3821), .Y(n3822) );
  INVX1 U4042 ( .A(n995), .Y(n3823) );
  INVX1 U4043 ( .A(n3823), .Y(n3824) );
  BUFX2 U4044 ( .A(n982), .Y(n3825) );
  INVX1 U4045 ( .A(n973), .Y(n3826) );
  INVX1 U4046 ( .A(n3826), .Y(n3827) );
  BUFX2 U4047 ( .A(n956), .Y(n3828) );
  INVX1 U4048 ( .A(n943), .Y(n3829) );
  INVX1 U4049 ( .A(n3829), .Y(n3830) );
  BUFX2 U4050 ( .A(n932), .Y(n3831) );
  INVX1 U4051 ( .A(n915), .Y(n3832) );
  INVX1 U4052 ( .A(n3832), .Y(n3833) );
  INVX1 U4053 ( .A(n904), .Y(n3834) );
  INVX1 U4054 ( .A(n3834), .Y(n3835) );
  INVX1 U4055 ( .A(n889), .Y(n3836) );
  INVX1 U4056 ( .A(n3836), .Y(n3837) );
  INVX1 U4057 ( .A(n878), .Y(n3838) );
  INVX1 U4058 ( .A(n3838), .Y(n3839) );
  INVX1 U4059 ( .A(n869), .Y(n3840) );
  INVX1 U4060 ( .A(n3840), .Y(n3841) );
  INVX1 U4061 ( .A(n861), .Y(n3842) );
  INVX1 U4062 ( .A(n3842), .Y(n3843) );
  BUFX2 U4063 ( .A(n824), .Y(n3844) );
  BUFX2 U4064 ( .A(n794), .Y(n3845) );
  BUFX2 U4065 ( .A(n777), .Y(n3846) );
  BUFX2 U4066 ( .A(n762), .Y(n3847) );
  BUFX2 U4067 ( .A(n749), .Y(n3848) );
  INVX1 U4068 ( .A(n745), .Y(n3849) );
  INVX1 U4069 ( .A(n3849), .Y(n3850) );
  INVX1 U4070 ( .A(n675), .Y(n3851) );
  INVX1 U4071 ( .A(n3851), .Y(n3852) );
  INVX1 U4072 ( .A(n593), .Y(n3853) );
  INVX1 U4073 ( .A(n3853), .Y(n3854) );
  INVX1 U4074 ( .A(n507), .Y(n3855) );
  INVX1 U4075 ( .A(n3855), .Y(n3856) );
  BUFX2 U4076 ( .A(n437), .Y(n3857) );
  INVX1 U4077 ( .A(n417), .Y(n3858) );
  INVX1 U4078 ( .A(n3858), .Y(n3859) );
  INVX1 U4079 ( .A(n331), .Y(n3860) );
  INVX1 U4080 ( .A(n3860), .Y(n3861) );
  BUFX2 U4081 ( .A(n261), .Y(n3862) );
  INVX1 U4082 ( .A(n241), .Y(n3863) );
  INVX1 U4083 ( .A(n3863), .Y(n3864) );
  BUFX2 U4084 ( .A(n208), .Y(n3865) );
  INVX1 U4085 ( .A(n4148), .Y(n3866) );
  INVX1 U4086 ( .A(n4759), .Y(n3867) );
  INVX1 U4087 ( .A(n4677), .Y(n3868) );
  INVX1 U4088 ( .A(n4720), .Y(n3869) );
  INVX1 U4089 ( .A(n3886), .Y(n3870) );
  INVX1 U4090 ( .A(n4480), .Y(n3871) );
  OR2X2 U4091 ( .A(n1765), .B(n4296), .Y(n1703) );
  INVX1 U4092 ( .A(n1703), .Y(n3872) );
  INVX1 U4093 ( .A(n1703), .Y(n3873) );
  INVX1 U4094 ( .A(n944), .Y(n3874) );
  AND2X2 U4095 ( .A(n2848), .B(n2929), .Y(n1226) );
  INVX1 U4096 ( .A(n1226), .Y(n3875) );
  INVX1 U4097 ( .A(n1226), .Y(n3876) );
  AND2X2 U4098 ( .A(n2848), .B(n2930), .Y(n1202) );
  INVX1 U4099 ( .A(n1202), .Y(n3877) );
  AND2X2 U4100 ( .A(n4597), .B(n584), .Y(n498) );
  INVX1 U4101 ( .A(n498), .Y(n3878) );
  INVX1 U4102 ( .A(n498), .Y(n3879) );
  INVX1 U4103 ( .A(n4768), .Y(n3880) );
  INVX1 U4104 ( .A(n1313), .Y(n3881) );
  INVX1 U4105 ( .A(n1289), .Y(n3882) );
  INVX1 U4106 ( .A(n1245), .Y(n3883) );
  INVX1 U4107 ( .A(n1225), .Y(n3884) );
  INVX1 U4108 ( .A(n2035), .Y(n3885) );
  INVX1 U4109 ( .A(n1846), .Y(n3887) );
  INVX1 U4110 ( .A(n1846), .Y(n3888) );
  INVX1 U4111 ( .A(n3435), .Y(n3889) );
  INVX1 U4112 ( .A(n464), .Y(n3890) );
  INVX1 U4113 ( .A(n4159), .Y(n3891) );
  INVX1 U4114 ( .A(n3893), .Y(n3892) );
  INVX1 U4115 ( .A(n3741), .Y(n3893) );
  INVX1 U4116 ( .A(n3743), .Y(n3894) );
  INVX1 U4117 ( .A(n3897), .Y(n3895) );
  INVX1 U4118 ( .A(n3895), .Y(n3896) );
  INVX1 U4119 ( .A(n3744), .Y(n3897) );
  INVX1 U4120 ( .A(n4345), .Y(n3898) );
  AND2X2 U4121 ( .A(B[179]), .B(A[179]), .Y(n199) );
  INVX1 U4122 ( .A(n199), .Y(n3899) );
  INVX1 U4123 ( .A(n4732), .Y(n3900) );
  INVX1 U4124 ( .A(n4173), .Y(n3901) );
  INVX1 U4125 ( .A(n4175), .Y(n3902) );
  INVX1 U4126 ( .A(n4185), .Y(n3903) );
  INVX1 U4127 ( .A(n4675), .Y(n3904) );
  INVX1 U4128 ( .A(n4666), .Y(n3905) );
  AND2X2 U4129 ( .A(n584), .B(n3116), .Y(n4159) );
  INVX1 U4130 ( .A(n4159), .Y(n3906) );
  INVX1 U4131 ( .A(n4493), .Y(n3907) );
  INVX1 U4132 ( .A(n4458), .Y(n3908) );
  INVX1 U4133 ( .A(n4713), .Y(n3909) );
  INVX1 U4134 ( .A(n4178), .Y(n3910) );
  INVX1 U4135 ( .A(n4497), .Y(n3911) );
  INVX1 U4136 ( .A(n4674), .Y(n3912) );
  INVX1 U4137 ( .A(n4706), .Y(n3913) );
  INVX1 U4138 ( .A(n4697), .Y(n3914) );
  INVX1 U4139 ( .A(n4676), .Y(n3915) );
  INVX1 U4140 ( .A(n4673), .Y(n3916) );
  INVX1 U4141 ( .A(n4663), .Y(n3917) );
  INVX1 U4142 ( .A(n1997), .Y(n3918) );
  OR2X2 U4143 ( .A(n1982), .B(n4780), .Y(n1975) );
  OR2X2 U4144 ( .A(n3398), .B(n4751), .Y(n1955) );
  INVX1 U4145 ( .A(n1955), .Y(n3919) );
  OR2X2 U4146 ( .A(n3181), .B(n4733), .Y(n1937) );
  INVX1 U4147 ( .A(n1937), .Y(n3920) );
  INVX1 U4148 ( .A(n1489), .Y(n3921) );
  OR2X2 U4149 ( .A(n1476), .B(n4765), .Y(n1467) );
  INVX1 U4150 ( .A(n1467), .Y(n3922) );
  OR2X2 U4151 ( .A(n4150), .B(n4442), .Y(n1429) );
  INVX1 U4152 ( .A(n1429), .Y(n3923) );
  OR2X2 U4153 ( .A(n4316), .B(n4756), .Y(n1405) );
  INVX1 U4154 ( .A(n1405), .Y(n3924) );
  OR2X2 U4155 ( .A(n3371), .B(n4766), .Y(n1387) );
  INVX1 U4156 ( .A(n1387), .Y(n3925) );
  OR2X2 U4157 ( .A(n4327), .B(n4435), .Y(n1365) );
  INVX1 U4158 ( .A(n1365), .Y(n3926) );
  OR2X2 U4159 ( .A(n3373), .B(n4664), .Y(n1347) );
  INVX1 U4160 ( .A(n1347), .Y(n3927) );
  OR2X2 U4161 ( .A(n3399), .B(n4431), .Y(n1323) );
  INVX1 U4162 ( .A(n1323), .Y(n3928) );
  OR2X2 U4163 ( .A(n3375), .B(n4433), .Y(n1305) );
  INVX1 U4164 ( .A(n1305), .Y(n3929) );
  OR2X2 U4165 ( .A(n3029), .B(n4412), .Y(n1281) );
  INVX1 U4166 ( .A(n1281), .Y(n3930) );
  OR2X2 U4167 ( .A(n3366), .B(n4428), .Y(n1261) );
  INVX1 U4168 ( .A(n1261), .Y(n3931) );
  OR2X2 U4169 ( .A(n3377), .B(n4408), .Y(n1237) );
  INVX1 U4170 ( .A(n1237), .Y(n3932) );
  INVX1 U4171 ( .A(n1086), .Y(n3933) );
  INVX1 U4172 ( .A(n875), .Y(n3934) );
  INVX1 U4173 ( .A(n858), .Y(n3935) );
  OR2X2 U4174 ( .A(n728), .B(n4420), .Y(n719) );
  INVX1 U4175 ( .A(n719), .Y(n3936) );
  OR2X2 U4176 ( .A(n4320), .B(n4470), .Y(n699) );
  INVX1 U4177 ( .A(n699), .Y(n3937) );
  OR2X2 U4178 ( .A(n3381), .B(n4397), .Y(n681) );
  INVX1 U4179 ( .A(n681), .Y(n3938) );
  OR2X2 U4180 ( .A(n670), .B(n4393), .Y(n657) );
  INVX1 U4181 ( .A(n657), .Y(n3939) );
  OR2X2 U4182 ( .A(n3383), .B(n4416), .Y(n639) );
  INVX1 U4183 ( .A(n639), .Y(n3940) );
  OR2X2 U4184 ( .A(n626), .B(n4386), .Y(n617) );
  INVX1 U4185 ( .A(n617), .Y(n3941) );
  OR2X2 U4186 ( .A(n3385), .B(n4374), .Y(n599) );
  INVX1 U4187 ( .A(n599), .Y(n3942) );
  OR2X2 U4188 ( .A(n4324), .B(n4604), .Y(n575) );
  INVX1 U4189 ( .A(n575), .Y(n3943) );
  OR2X2 U4190 ( .A(n3387), .B(n4372), .Y(n557) );
  INVX1 U4191 ( .A(n557), .Y(n3944) );
  OR2X2 U4192 ( .A(n3389), .B(n4608), .Y(n533) );
  INVX1 U4193 ( .A(n533), .Y(n3945) );
  OR2X2 U4194 ( .A(n3391), .B(n4369), .Y(n513) );
  INVX1 U4195 ( .A(n513), .Y(n3946) );
  OR2X2 U4196 ( .A(n3878), .B(n4610), .Y(n489) );
  INVX1 U4197 ( .A(n489), .Y(n3947) );
  OR2X2 U4198 ( .A(n3906), .B(n4612), .Y(n469) );
  INVX1 U4199 ( .A(n469), .Y(n3948) );
  OR2X2 U4200 ( .A(n4160), .B(n4613), .Y(n423) );
  INVX1 U4201 ( .A(n423), .Y(n3949) );
  AND2X2 U4202 ( .A(n2048), .B(n3731), .Y(n2044) );
  INVX1 U4203 ( .A(n2044), .Y(n3950) );
  AND2X2 U4204 ( .A(n2275), .B(n2035), .Y(n2026) );
  INVX1 U4205 ( .A(n2026), .Y(n3951) );
  AND2X2 U4206 ( .A(n4763), .B(n2035), .Y(n2015) );
  INVX1 U4207 ( .A(n2015), .Y(n3952) );
  AND2X2 U4208 ( .A(n2035), .B(n4257), .Y(n2006) );
  INVX1 U4209 ( .A(n2006), .Y(n3953) );
  AND2X2 U4210 ( .A(n2253), .B(n4314), .Y(n1816) );
  INVX1 U4211 ( .A(n1816), .Y(n3954) );
  AND2X2 U4212 ( .A(n2251), .B(n1803), .Y(n1794) );
  INVX1 U4213 ( .A(n1794), .Y(n3955) );
  AND2X2 U4214 ( .A(n2891), .B(n3271), .Y(n1776) );
  INVX1 U4215 ( .A(n1776), .Y(n3956) );
  AND2X2 U4216 ( .A(n1758), .B(n4315), .Y(n1754) );
  INVX1 U4217 ( .A(n1754), .Y(n3957) );
  AND2X2 U4218 ( .A(n1740), .B(n4133), .Y(n1736) );
  INVX1 U4219 ( .A(n1736), .Y(n3958) );
  AND2X2 U4220 ( .A(n4170), .B(n4135), .Y(n1714) );
  INVX1 U4221 ( .A(n1714), .Y(n3959) );
  AND2X2 U4222 ( .A(n4149), .B(n3872), .Y(n1694) );
  INVX1 U4223 ( .A(n1694), .Y(n3960) );
  AND2X2 U4224 ( .A(n1676), .B(n1681), .Y(n1672) );
  INVX1 U4225 ( .A(n1672), .Y(n3961) );
  AND2X2 U4226 ( .A(n4592), .B(n1681), .Y(n1661) );
  INVX1 U4227 ( .A(n1661), .Y(n3962) );
  AND2X2 U4228 ( .A(n4276), .B(n1681), .Y(n1652) );
  INVX1 U4229 ( .A(n1652), .Y(n3963) );
  AND2X2 U4230 ( .A(n2861), .B(n1681), .Y(n1637) );
  INVX1 U4231 ( .A(n1637), .Y(n3964) );
  AND2X2 U4232 ( .A(n2925), .B(n1681), .Y(n1628) );
  INVX1 U4233 ( .A(n1628), .Y(n3965) );
  AND2X2 U4234 ( .A(n1617), .B(n1681), .Y(n1615) );
  INVX1 U4235 ( .A(n1615), .Y(n3966) );
  AND2X2 U4236 ( .A(n2926), .B(n1681), .Y(n1606) );
  INVX1 U4237 ( .A(n1606), .Y(n3967) );
  INVX1 U4238 ( .A(n1591), .Y(n3968) );
  AND2X2 U4239 ( .A(n4739), .B(n1681), .Y(n1591) );
  AND2X2 U4240 ( .A(n1681), .B(n3007), .Y(n1582) );
  INVX1 U4241 ( .A(n1582), .Y(n3969) );
  AND2X2 U4242 ( .A(n1681), .B(n3009), .Y(n1567) );
  INVX1 U4243 ( .A(n1567), .Y(n3970) );
  AND2X2 U4244 ( .A(n1681), .B(n3010), .Y(n1556) );
  INVX1 U4245 ( .A(n1556), .Y(n3971) );
  AND2X2 U4246 ( .A(n1681), .B(n3012), .Y(n1541) );
  INVX1 U4247 ( .A(n1541), .Y(n3972) );
  AND2X2 U4248 ( .A(n1681), .B(n3013), .Y(n1530) );
  INVX1 U4249 ( .A(n1530), .Y(n3973) );
  AND2X2 U4250 ( .A(n1681), .B(n3016), .Y(n1515) );
  INVX1 U4251 ( .A(n1515), .Y(n3974) );
  AND2X2 U4252 ( .A(n1681), .B(n2901), .Y(n1502) );
  INVX1 U4253 ( .A(n1502), .Y(n3975) );
  INVX1 U4254 ( .A(n2130), .Y(n3976) );
  INVX1 U4255 ( .A(n3978), .Y(n3977) );
  INVX1 U4256 ( .A(n4497), .Y(n3978) );
  INVX1 U4257 ( .A(n2023), .Y(n3979) );
  BUFX2 U4258 ( .A(n1848), .Y(n3980) );
  AND2X2 U4259 ( .A(n2957), .B(n2870), .Y(n194) );
  AND2X2 U4260 ( .A(n2962), .B(n4754), .Y(n188) );
  INVX1 U4261 ( .A(n188), .Y(n3981) );
  AND2X2 U4262 ( .A(n2963), .B(n2905), .Y(n186) );
  INVX1 U4263 ( .A(n186), .Y(n3982) );
  AND2X2 U4264 ( .A(n3208), .B(n2275), .Y(n185) );
  INVX1 U4265 ( .A(n185), .Y(n3983) );
  AND2X2 U4266 ( .A(n4190), .B(n2023), .Y(n184) );
  INVX1 U4267 ( .A(n184), .Y(n3984) );
  AND2X2 U4268 ( .A(n3511), .B(n4402), .Y(n183) );
  INVX1 U4269 ( .A(n183), .Y(n3985) );
  AND2X2 U4270 ( .A(n4191), .B(n4448), .Y(n182) );
  INVX1 U4271 ( .A(n182), .Y(n3986) );
  AND2X2 U4272 ( .A(n3894), .B(n1993), .Y(n181) );
  AND2X2 U4273 ( .A(n3288), .B(n4768), .Y(n164) );
  INVX1 U4274 ( .A(n164), .Y(n3987) );
  AND2X2 U4275 ( .A(n4646), .B(n2253), .Y(n163) );
  INVX1 U4276 ( .A(n163), .Y(n3988) );
  AND2X2 U4277 ( .A(n2989), .B(n1813), .Y(n162) );
  INVX1 U4278 ( .A(n162), .Y(n3989) );
  AND2X2 U4279 ( .A(n4344), .B(n2251), .Y(n161) );
  INVX1 U4280 ( .A(n161), .Y(n3990) );
  AND2X2 U4281 ( .A(n4193), .B(n2250), .Y(n160) );
  INVX1 U4282 ( .A(n160), .Y(n3991) );
  AND2X2 U4283 ( .A(n2991), .B(n2891), .Y(n159) );
  INVX1 U4284 ( .A(n159), .Y(n3992) );
  AND2X2 U4285 ( .A(n2992), .B(n2248), .Y(n158) );
  INVX1 U4286 ( .A(n158), .Y(n3993) );
  AND2X2 U4287 ( .A(n3223), .B(n1758), .Y(n157) );
  INVX1 U4288 ( .A(n157), .Y(n3994) );
  AND2X2 U4289 ( .A(n2994), .B(n4477), .Y(n156) );
  INVX1 U4290 ( .A(n156), .Y(n3995) );
  AND2X2 U4291 ( .A(n3499), .B(n1740), .Y(n155) );
  INVX1 U4292 ( .A(n155), .Y(n3996) );
  AND2X2 U4293 ( .A(n2995), .B(n2244), .Y(n154) );
  INVX1 U4294 ( .A(n154), .Y(n3997) );
  AND2X2 U4295 ( .A(n2998), .B(n2242), .Y(n152) );
  INVX1 U4296 ( .A(n152), .Y(n3998) );
  AND2X2 U4297 ( .A(n4356), .B(n4149), .Y(n151) );
  INVX1 U4298 ( .A(n151), .Y(n3999) );
  AND2X2 U4299 ( .A(n3000), .B(n2240), .Y(n150) );
  INVX1 U4300 ( .A(n150), .Y(n4000) );
  AND2X2 U4301 ( .A(n3896), .B(n1676), .Y(n149) );
  INVX1 U4302 ( .A(n149), .Y(n4001) );
  AND2X2 U4303 ( .A(n3001), .B(n3886), .Y(n148) );
  INVX1 U4304 ( .A(n148), .Y(n4002) );
  AND2X2 U4305 ( .A(n4551), .B(n1656), .Y(n147) );
  AND2X2 U4306 ( .A(n3002), .B(n2236), .Y(n146) );
  INVX1 U4307 ( .A(n146), .Y(n4003) );
  AND2X2 U4308 ( .A(n3003), .B(n4480), .Y(n144) );
  INVX1 U4309 ( .A(n144), .Y(n4004) );
  AND2X2 U4310 ( .A(n2919), .B(n2233), .Y(n143) );
  INVX1 U4311 ( .A(n143), .Y(n4005) );
  AND2X2 U4312 ( .A(n3004), .B(n2232), .Y(n142) );
  INVX1 U4313 ( .A(n142), .Y(n4006) );
  AND2X2 U4314 ( .A(n2920), .B(n2231), .Y(n141) );
  INVX1 U4315 ( .A(n141), .Y(n4007) );
  AND2X2 U4316 ( .A(n3008), .B(n1579), .Y(n140) );
  INVX1 U4317 ( .A(n140), .Y(n4008) );
  AND2X2 U4318 ( .A(n3211), .B(n2229), .Y(n139) );
  INVX1 U4319 ( .A(n139), .Y(n4009) );
  AND2X2 U4320 ( .A(n3011), .B(n2228), .Y(n138) );
  INVX1 U4321 ( .A(n138), .Y(n4010) );
  AND2X2 U4322 ( .A(n3212), .B(n2227), .Y(n137) );
  INVX1 U4323 ( .A(n137), .Y(n4011) );
  AND2X2 U4324 ( .A(n3014), .B(n2226), .Y(n136) );
  INVX1 U4325 ( .A(n136), .Y(n4012) );
  AND2X2 U4326 ( .A(n4552), .B(n2225), .Y(n135) );
  INVX1 U4327 ( .A(n135), .Y(n4013) );
  AND2X2 U4328 ( .A(n3018), .B(n2224), .Y(n134) );
  INVX1 U4329 ( .A(n134), .Y(n4014) );
  AND2X2 U4330 ( .A(n3473), .B(n1485), .Y(n133) );
  AND2X2 U4331 ( .A(n4354), .B(n737), .Y(n69) );
  INVX1 U4332 ( .A(n69), .Y(n4015) );
  AND2X2 U4333 ( .A(n2959), .B(n4694), .Y(n191) );
  INVX1 U4334 ( .A(n191), .Y(n4016) );
  AND2X2 U4335 ( .A(n2965), .B(n2270), .Y(n180) );
  INVX1 U4336 ( .A(n180), .Y(n4017) );
  AND2X2 U4337 ( .A(n2967), .B(n2268), .Y(n178) );
  INVX1 U4338 ( .A(n178), .Y(n4018) );
  AND2X2 U4339 ( .A(n2915), .B(n4144), .Y(n177) );
  INVX1 U4340 ( .A(n177), .Y(n4019) );
  AND2X2 U4341 ( .A(n2969), .B(n2266), .Y(n176) );
  INVX1 U4342 ( .A(n176), .Y(n4020) );
  AND2X2 U4343 ( .A(n4192), .B(n2264), .Y(n174) );
  INVX1 U4344 ( .A(n174), .Y(n4021) );
  AND2X2 U4345 ( .A(n3209), .B(n1919), .Y(n173) );
  INVX1 U4346 ( .A(n173), .Y(n4022) );
  AND2X2 U4347 ( .A(n3210), .B(n4148), .Y(n169) );
  INVX1 U4348 ( .A(n169), .Y(n4023) );
  AND2X2 U4349 ( .A(n2981), .B(n2258), .Y(n168) );
  INVX1 U4350 ( .A(n168), .Y(n4024) );
  AND2X2 U4351 ( .A(n2985), .B(n4422), .Y(n167) );
  INVX1 U4352 ( .A(n167), .Y(n4025) );
  AND2X2 U4353 ( .A(n2987), .B(n1846), .Y(n166) );
  INVX1 U4354 ( .A(n166), .Y(n4026) );
  AND2X2 U4355 ( .A(n3513), .B(n1834), .Y(n165) );
  AND2X2 U4356 ( .A(n3019), .B(n2222), .Y(n132) );
  INVX1 U4357 ( .A(n132), .Y(n4027) );
  AND2X2 U4358 ( .A(n2921), .B(n2221), .Y(n131) );
  INVX1 U4359 ( .A(n131), .Y(n4028) );
  AND2X2 U4360 ( .A(n3020), .B(n4174), .Y(n130) );
  INVX1 U4361 ( .A(n130), .Y(n4029) );
  AND2X2 U4362 ( .A(n2916), .B(n4444), .Y(n129) );
  INVX1 U4363 ( .A(n129), .Y(n4030) );
  AND2X2 U4364 ( .A(n4194), .B(n2218), .Y(n128) );
  INVX1 U4365 ( .A(n128), .Y(n4031) );
  AND2X2 U4366 ( .A(n3507), .B(n4440), .Y(n127) );
  INVX1 U4367 ( .A(n127), .Y(n4032) );
  AND2X2 U4368 ( .A(n4195), .B(n2216), .Y(n126) );
  INVX1 U4369 ( .A(n126), .Y(n4033) );
  AND2X2 U4370 ( .A(n3219), .B(n4175), .Y(n125) );
  INVX1 U4371 ( .A(n125), .Y(n4034) );
  AND2X2 U4372 ( .A(n3022), .B(n2214), .Y(n124) );
  INVX1 U4373 ( .A(n124), .Y(n4035) );
  AND2X2 U4374 ( .A(n2922), .B(n1389), .Y(n123) );
  INVX1 U4375 ( .A(n123), .Y(n4036) );
  AND2X2 U4376 ( .A(n3024), .B(n1384), .Y(n122) );
  INVX1 U4377 ( .A(n122), .Y(n4037) );
  AND2X2 U4378 ( .A(n4554), .B(n2211), .Y(n121) );
  INVX1 U4379 ( .A(n121), .Y(n4038) );
  AND2X2 U4380 ( .A(n3026), .B(n4176), .Y(n120) );
  INVX1 U4381 ( .A(n120), .Y(n4039) );
  AND2X2 U4382 ( .A(n3027), .B(n4771), .Y(n119) );
  INVX1 U4383 ( .A(n119), .Y(n4040) );
  AND2X2 U4384 ( .A(n4196), .B(n2208), .Y(n118) );
  INVX1 U4385 ( .A(n118), .Y(n4041) );
  AND2X2 U4386 ( .A(n3475), .B(n2207), .Y(n117) );
  INVX1 U4387 ( .A(n117), .Y(n4042) );
  AND2X2 U4388 ( .A(n4197), .B(n1320), .Y(n116) );
  INVX1 U4389 ( .A(n116), .Y(n4043) );
  AND2X2 U4390 ( .A(n2928), .B(n2205), .Y(n115) );
  INVX1 U4391 ( .A(n115), .Y(n4044) );
  AND2X2 U4392 ( .A(n4198), .B(n2204), .Y(n114) );
  INVX1 U4393 ( .A(n114), .Y(n4045) );
  AND2X2 U4394 ( .A(n3030), .B(n2203), .Y(n113) );
  INVX1 U4395 ( .A(n113), .Y(n4046) );
  AND2X2 U4396 ( .A(n4199), .B(n2202), .Y(n112) );
  INVX1 U4397 ( .A(n112), .Y(n4047) );
  AND2X2 U4398 ( .A(n4556), .B(n4426), .Y(n111) );
  INVX1 U4399 ( .A(n111), .Y(n4048) );
  AND2X2 U4400 ( .A(n4200), .B(n2200), .Y(n110) );
  INVX1 U4401 ( .A(n110), .Y(n4049) );
  AND2X2 U4402 ( .A(n4557), .B(n2199), .Y(n109) );
  INVX1 U4403 ( .A(n109), .Y(n4050) );
  AND2X2 U4404 ( .A(n4201), .B(n1234), .Y(n108) );
  INVX1 U4405 ( .A(n108), .Y(n4051) );
  AND2X2 U4406 ( .A(n3033), .B(n1219), .Y(n107) );
  INVX1 U4407 ( .A(n107), .Y(n4052) );
  AND2X2 U4408 ( .A(n3035), .B(n4178), .Y(n106) );
  INVX1 U4409 ( .A(n106), .Y(n4053) );
  AND2X2 U4410 ( .A(n2931), .B(n2195), .Y(n105) );
  INVX1 U4411 ( .A(n105), .Y(n4054) );
  AND2X2 U4412 ( .A(n4202), .B(n4166), .Y(n104) );
  INVX1 U4413 ( .A(n104), .Y(n4055) );
  AND2X2 U4414 ( .A(n2955), .B(n4759), .Y(n103) );
  INVX1 U4415 ( .A(n103), .Y(n4056) );
  AND2X2 U4416 ( .A(n3039), .B(n1168), .Y(n102) );
  INVX1 U4417 ( .A(n102), .Y(n4057) );
  AND2X2 U4418 ( .A(n3220), .B(n2191), .Y(n101) );
  INVX1 U4419 ( .A(n101), .Y(n4058) );
  AND2X2 U4420 ( .A(n3042), .B(n4247), .Y(n100) );
  INVX1 U4421 ( .A(n100), .Y(n4059) );
  AND2X2 U4422 ( .A(n3045), .B(n2188), .Y(n98) );
  INVX1 U4423 ( .A(n98), .Y(n4060) );
  AND2X2 U4424 ( .A(n3898), .B(n2187), .Y(n97) );
  INVX1 U4425 ( .A(n97), .Y(n4061) );
  AND2X2 U4426 ( .A(n3049), .B(n3907), .Y(n96) );
  INVX1 U4427 ( .A(n96), .Y(n4062) );
  AND2X2 U4428 ( .A(n4347), .B(n4181), .Y(n95) );
  INVX1 U4429 ( .A(n95), .Y(n4063) );
  AND2X2 U4430 ( .A(n3050), .B(n2184), .Y(n94) );
  INVX1 U4431 ( .A(n94), .Y(n4064) );
  AND2X2 U4432 ( .A(n3213), .B(n3752), .Y(n93) );
  INVX1 U4433 ( .A(n93), .Y(n4065) );
  AND2X2 U4434 ( .A(n4203), .B(n2182), .Y(n92) );
  INVX1 U4435 ( .A(n92), .Y(n4066) );
  AND2X2 U4436 ( .A(n4348), .B(n2181), .Y(n91) );
  INVX1 U4437 ( .A(n91), .Y(n4067) );
  AND2X2 U4438 ( .A(n3058), .B(n2180), .Y(n90) );
  INVX1 U4439 ( .A(n90), .Y(n4068) );
  AND2X2 U4440 ( .A(n4349), .B(n1009), .Y(n89) );
  INVX1 U4441 ( .A(n89), .Y(n4069) );
  AND2X2 U4442 ( .A(n3063), .B(n3977), .Y(n88) );
  INVX1 U4443 ( .A(n88), .Y(n4070) );
  AND2X2 U4444 ( .A(n4351), .B(n4184), .Y(n87) );
  INVX1 U4445 ( .A(n87), .Y(n4071) );
  AND2X2 U4446 ( .A(n3067), .B(n2176), .Y(n86) );
  INVX1 U4447 ( .A(n86), .Y(n4072) );
  AND2X2 U4448 ( .A(n3214), .B(n959), .Y(n85) );
  INVX1 U4449 ( .A(n85), .Y(n4073) );
  AND2X2 U4450 ( .A(n3072), .B(n3889), .Y(n84) );
  INVX1 U4451 ( .A(n84), .Y(n4074) );
  AND2X2 U4452 ( .A(n4558), .B(n2173), .Y(n83) );
  INVX1 U4453 ( .A(n83), .Y(n4075) );
  AND2X2 U4454 ( .A(n3075), .B(n926), .Y(n82) );
  INVX1 U4455 ( .A(n82), .Y(n4076) );
  AND2X2 U4456 ( .A(n3479), .B(n4376), .Y(n81) );
  INVX1 U4457 ( .A(n81), .Y(n4077) );
  AND2X2 U4458 ( .A(n3076), .B(n898), .Y(n80) );
  INVX1 U4459 ( .A(n80), .Y(n4078) );
  AND2X2 U4460 ( .A(n4559), .B(n4388), .Y(n79) );
  INVX1 U4461 ( .A(n79), .Y(n4079) );
  AND2X2 U4462 ( .A(n3079), .B(n4185), .Y(n78) );
  INVX1 U4463 ( .A(n78), .Y(n4080) );
  AND2X2 U4464 ( .A(n4560), .B(n2167), .Y(n77) );
  INVX1 U4465 ( .A(n77), .Y(n4081) );
  AND2X2 U4466 ( .A(n3083), .B(n2166), .Y(n76) );
  INVX1 U4467 ( .A(n76), .Y(n4082) );
  AND2X2 U4468 ( .A(n4352), .B(n827), .Y(n75) );
  INVX1 U4469 ( .A(n75), .Y(n4083) );
  AND2X2 U4470 ( .A(n3084), .B(n2164), .Y(n74) );
  INVX1 U4471 ( .A(n74), .Y(n4084) );
  AND2X2 U4472 ( .A(n3215), .B(n795), .Y(n73) );
  INVX1 U4473 ( .A(n73), .Y(n4085) );
  AND2X2 U4474 ( .A(n3087), .B(n784), .Y(n72) );
  INVX1 U4475 ( .A(n72), .Y(n4086) );
  AND2X2 U4476 ( .A(n4561), .B(n4380), .Y(n71) );
  INVX1 U4477 ( .A(n71), .Y(n4087) );
  AND2X2 U4478 ( .A(n3090), .B(n2160), .Y(n70) );
  INVX1 U4479 ( .A(n70), .Y(n4088) );
  AND2X2 U4480 ( .A(n4204), .B(n2158), .Y(n68) );
  INVX1 U4481 ( .A(n68), .Y(n4089) );
  AND2X2 U4482 ( .A(n3471), .B(n4418), .Y(n67) );
  INVX1 U4483 ( .A(n67), .Y(n4090) );
  AND2X2 U4484 ( .A(n3093), .B(n2156), .Y(n66) );
  INVX1 U4485 ( .A(n66), .Y(n4091) );
  AND2X2 U4486 ( .A(n2917), .B(n2155), .Y(n65) );
  INVX1 U4487 ( .A(n65), .Y(n4092) );
  AND2X2 U4488 ( .A(n3095), .B(n4250), .Y(n64) );
  INVX1 U4489 ( .A(n64), .Y(n4093) );
  AND2X2 U4490 ( .A(n2923), .B(n4395), .Y(n63) );
  INVX1 U4491 ( .A(n63), .Y(n4094) );
  AND2X2 U4492 ( .A(n3096), .B(n2152), .Y(n62) );
  INVX1 U4493 ( .A(n62), .Y(n4095) );
  AND2X2 U4494 ( .A(n4562), .B(n2151), .Y(n61) );
  INVX1 U4495 ( .A(n61), .Y(n4096) );
  AND2X2 U4496 ( .A(n3099), .B(n654), .Y(n60) );
  INVX1 U4497 ( .A(n60), .Y(n4097) );
  AND2X2 U4498 ( .A(n4563), .B(n2149), .Y(n59) );
  INVX1 U4499 ( .A(n59), .Y(n4098) );
  AND2X2 U4500 ( .A(n3100), .B(n2148), .Y(n58) );
  INVX1 U4501 ( .A(n58), .Y(n4099) );
  AND2X2 U4502 ( .A(n3485), .B(n4384), .Y(n57) );
  INVX1 U4503 ( .A(n57), .Y(n4100) );
  AND2X2 U4504 ( .A(n3104), .B(n614), .Y(n56) );
  INVX1 U4505 ( .A(n56), .Y(n4101) );
  AND2X2 U4506 ( .A(n3106), .B(n2144), .Y(n54) );
  INVX1 U4507 ( .A(n54), .Y(n4102) );
  AND2X2 U4508 ( .A(n4565), .B(n2143), .Y(n53) );
  INVX1 U4509 ( .A(n53), .Y(n4103) );
  AND2X2 U4510 ( .A(n4205), .B(n572), .Y(n52) );
  INVX1 U4511 ( .A(n52), .Y(n4104) );
  AND2X2 U4512 ( .A(n2942), .B(n4670), .Y(n51) );
  INVX1 U4513 ( .A(n51), .Y(n4105) );
  AND2X2 U4514 ( .A(n4206), .B(n2140), .Y(n50) );
  INVX1 U4515 ( .A(n50), .Y(n4106) );
  AND2X2 U4516 ( .A(n4207), .B(n2138), .Y(n48) );
  INVX1 U4517 ( .A(n48), .Y(n4107) );
  AND2X2 U4518 ( .A(n4208), .B(n2136), .Y(n46) );
  INVX1 U4519 ( .A(n46), .Y(n4108) );
  AND2X2 U4520 ( .A(n4567), .B(n2135), .Y(n45) );
  INVX1 U4521 ( .A(n45), .Y(n4109) );
  AND2X2 U4522 ( .A(n3114), .B(n2134), .Y(n44) );
  INVX1 U4523 ( .A(n44), .Y(n4110) );
  AND2X2 U4524 ( .A(n4569), .B(n2133), .Y(n43) );
  INVX1 U4525 ( .A(n43), .Y(n4111) );
  AND2X2 U4526 ( .A(n4571), .B(n4364), .Y(n41) );
  INVX1 U4527 ( .A(n41), .Y(n4112) );
  AND2X2 U4528 ( .A(n3119), .B(n2130), .Y(n40) );
  INVX1 U4529 ( .A(n40), .Y(n4113) );
  AND2X2 U4530 ( .A(n4573), .B(n2129), .Y(n39) );
  INVX1 U4531 ( .A(n39), .Y(n4114) );
  AND2X2 U4532 ( .A(n3122), .B(n2128), .Y(n38) );
  INVX1 U4533 ( .A(n38), .Y(n4115) );
  AND2X2 U4534 ( .A(n4575), .B(n2127), .Y(n37) );
  INVX1 U4535 ( .A(n37), .Y(n4116) );
  AND2X2 U4536 ( .A(n4209), .B(n2126), .Y(n36) );
  INVX1 U4537 ( .A(n36), .Y(n4117) );
  AND2X2 U4538 ( .A(n3489), .B(n2125), .Y(n35) );
  INVX1 U4539 ( .A(n35), .Y(n4118) );
  AND2X2 U4540 ( .A(n3217), .B(n2123), .Y(n33) );
  INVX1 U4541 ( .A(n33), .Y(n4119) );
  AND2X2 U4542 ( .A(n3129), .B(n354), .Y(n32) );
  INVX1 U4543 ( .A(n32), .Y(n4120) );
  AND2X2 U4544 ( .A(n3131), .B(n2120), .Y(n30) );
  INVX1 U4545 ( .A(n30), .Y(n4121) );
  AND2X2 U4546 ( .A(n3134), .B(n2118), .Y(n28) );
  INVX1 U4547 ( .A(n28), .Y(n4122) );
  AND2X2 U4548 ( .A(n4576), .B(n2117), .Y(n27) );
  INVX1 U4549 ( .A(n27), .Y(n4123) );
  AND2X2 U4550 ( .A(n3136), .B(n290), .Y(n26) );
  INVX1 U4551 ( .A(n26), .Y(n4124) );
  AND2X2 U4552 ( .A(n3523), .B(n2115), .Y(n25) );
  INVX1 U4553 ( .A(n25), .Y(n4125) );
  AND2X2 U4554 ( .A(n3365), .B(n2114), .Y(n24) );
  INVX1 U4555 ( .A(n24), .Y(n4126) );
  AND2X2 U4556 ( .A(n4577), .B(n2113), .Y(n23) );
  INVX1 U4557 ( .A(n23), .Y(n4127) );
  AND2X2 U4558 ( .A(n3140), .B(n244), .Y(n22) );
  INVX1 U4559 ( .A(n22), .Y(n4128) );
  AND2X2 U4560 ( .A(n3493), .B(n2111), .Y(n21) );
  INVX1 U4561 ( .A(n21), .Y(n4129) );
  AND2X2 U4562 ( .A(n3143), .B(n220), .Y(n20) );
  INVX1 U4563 ( .A(n20), .Y(n4130) );
  AND2X2 U4564 ( .A(n4143), .B(n4783), .Y(n19) );
  INVX1 U4565 ( .A(n19), .Y(n4131) );
  AND2X2 U4566 ( .A(n3899), .B(n4785), .Y(n18) );
  INVX1 U4567 ( .A(n18), .Y(n4132) );
  OR2X2 U4568 ( .A(n1765), .B(n1747), .Y(n1745) );
  INVX1 U4569 ( .A(n1745), .Y(n4133) );
  INVX1 U4570 ( .A(n1745), .Y(n4134) );
  OR2X2 U4571 ( .A(n1765), .B(n4699), .Y(n1723) );
  INVX1 U4572 ( .A(n1723), .Y(n4135) );
  INVX1 U4573 ( .A(n1723), .Y(n4136) );
  OR2X2 U4574 ( .A(n1064), .B(n1044), .Y(n1042) );
  INVX1 U4575 ( .A(n1042), .Y(n4137) );
  INVX1 U4576 ( .A(n1647), .Y(n4139) );
  INVX1 U4577 ( .A(n1493), .Y(n4140) );
  INVX1 U4578 ( .A(n1338), .Y(n4141) );
  AND2X2 U4579 ( .A(B[178]), .B(A[178]), .Y(n212) );
  INVX1 U4580 ( .A(n212), .Y(n4142) );
  INVX1 U4581 ( .A(n212), .Y(n4143) );
  INVX1 U4582 ( .A(n1919), .Y(n4147) );
  AND2X2 U4583 ( .A(n3300), .B(n4714), .Y(n1438) );
  INVX1 U4584 ( .A(n1438), .Y(n4150) );
  INVX1 U4585 ( .A(n1438), .Y(n4151) );
  INVX1 U4586 ( .A(n1234), .Y(n4153) );
  INVX1 U4587 ( .A(n1219), .Y(n4154) );
  AND2X2 U4588 ( .A(n2848), .B(n2932), .Y(n1180) );
  INVX1 U4589 ( .A(n1180), .Y(n4155) );
  INVX1 U4590 ( .A(n1180), .Y(n4156) );
  INVX1 U4591 ( .A(n926), .Y(n4157) );
  INVX1 U4592 ( .A(n737), .Y(n4158) );
  AND2X2 U4593 ( .A(n584), .B(n3121), .Y(n432) );
  INVX1 U4594 ( .A(n432), .Y(n4160) );
  INVX1 U4595 ( .A(n432), .Y(n4161) );
  INVX1 U4596 ( .A(n354), .Y(n4162) );
  INVX1 U4597 ( .A(n220), .Y(n4164) );
  AND2X2 U4598 ( .A(B[155]), .B(A[155]), .Y(n467) );
  INVX1 U4599 ( .A(n467), .Y(n4165) );
  INVX1 U4600 ( .A(n2023), .Y(n4167) );
  INVX1 U4601 ( .A(n1632), .Y(n4172) );
  INVX1 U4602 ( .A(n1258), .Y(n4177) );
  INVX1 U4603 ( .A(n572), .Y(n4187) );
  INVX1 U4604 ( .A(n290), .Y(n4188) );
  INVX1 U4605 ( .A(n244), .Y(n4189) );
  AND2X2 U4606 ( .A(B[13]), .B(A[13]), .Y(n2024) );
  INVX1 U4607 ( .A(n2024), .Y(n4190) );
  AND2X2 U4608 ( .A(B[15]), .B(A[15]), .Y(n2004) );
  INVX1 U4609 ( .A(n2004), .Y(n4191) );
  AND2X2 U4610 ( .A(B[23]), .B(A[23]), .Y(n1935) );
  INVX1 U4611 ( .A(n1935), .Y(n4192) );
  AND2X2 U4612 ( .A(B[37]), .B(A[37]), .Y(n1792) );
  INVX1 U4613 ( .A(n1792), .Y(n4193) );
  AND2X2 U4614 ( .A(B[69]), .B(A[69]), .Y(n1445) );
  INVX1 U4615 ( .A(n1445), .Y(n4194) );
  AND2X2 U4616 ( .A(B[71]), .B(A[71]), .Y(n1427) );
  INVX1 U4617 ( .A(n1427), .Y(n4195) );
  AND2X2 U4618 ( .A(B[79]), .B(A[79]), .Y(n1345) );
  INVX1 U4619 ( .A(n1345), .Y(n4196) );
  AND2X2 U4620 ( .A(B[81]), .B(A[81]), .Y(n1321) );
  INVX1 U4621 ( .A(n1321), .Y(n4197) );
  AND2X2 U4622 ( .A(B[83]), .B(A[83]), .Y(n1303) );
  INVX1 U4623 ( .A(n1303), .Y(n4198) );
  AND2X2 U4624 ( .A(B[85]), .B(A[85]), .Y(n1279) );
  INVX1 U4625 ( .A(n1279), .Y(n4199) );
  AND2X2 U4626 ( .A(B[87]), .B(A[87]), .Y(n1259) );
  INVX1 U4627 ( .A(n1259), .Y(n4200) );
  AND2X2 U4628 ( .A(B[89]), .B(A[89]), .Y(n1235) );
  INVX1 U4629 ( .A(n1235), .Y(n4201) );
  AND2X2 U4630 ( .A(B[93]), .B(A[93]), .Y(n1191) );
  INVX1 U4631 ( .A(n1191), .Y(n4202) );
  AND2X2 U4632 ( .A(B[105]), .B(A[105]), .Y(n1049) );
  INVX1 U4633 ( .A(n1049), .Y(n4203) );
  AND2X2 U4634 ( .A(B[129]), .B(A[129]), .Y(n733) );
  INVX1 U4635 ( .A(n733), .Y(n4204) );
  AND2X2 U4636 ( .A(B[145]), .B(A[145]), .Y(n573) );
  INVX1 U4637 ( .A(n573), .Y(n4205) );
  AND2X2 U4638 ( .A(B[147]), .B(A[147]), .Y(n555) );
  INVX1 U4639 ( .A(n555), .Y(n4206) );
  AND2X2 U4640 ( .A(B[149]), .B(A[149]), .Y(n531) );
  INVX1 U4641 ( .A(n531), .Y(n4207) );
  AND2X2 U4642 ( .A(B[151]), .B(A[151]), .Y(n511) );
  INVX1 U4643 ( .A(n511), .Y(n4208) );
  AND2X2 U4644 ( .A(B[161]), .B(A[161]), .Y(n397) );
  INVX1 U4645 ( .A(n397), .Y(n4209) );
  INVX1 U4646 ( .A(n1970), .Y(n4210) );
  INVX1 U4647 ( .A(n1168), .Y(n4216) );
  INVX1 U4648 ( .A(n1422), .Y(n4217) );
  INVX1 U4649 ( .A(n298), .Y(n4218) );
  INVX1 U4650 ( .A(n252), .Y(n4219) );
  INVX1 U4651 ( .A(n1945), .Y(n4230) );
  INVX1 U4652 ( .A(n1618), .Y(n4231) );
  INVX1 U4653 ( .A(n1437), .Y(n4232) );
  INVX1 U4654 ( .A(n1269), .Y(n4233) );
  INVX1 U4655 ( .A(n1201), .Y(n4234) );
  AOI21X1 U4656 ( .A(n1335), .B(n2932), .C(n1183), .Y(n4235) );
  INVX1 U4657 ( .A(n891), .Y(n4236) );
  INVX1 U4658 ( .A(n689), .Y(n4237) );
  INVX1 U4659 ( .A(n565), .Y(n4238) );
  INVX1 U4660 ( .A(n541), .Y(n4239) );
  INVX1 U4661 ( .A(n521), .Y(n4240) );
  INVX1 U4662 ( .A(n497), .Y(n4241) );
  INVX1 U4663 ( .A(n1513), .Y(n4243) );
  INVX1 U4664 ( .A(n1352), .Y(n4244) );
  INVX1 U4665 ( .A(n1222), .Y(n4245) );
  INVX1 U4666 ( .A(n4331), .Y(n4246) );
  INVX1 U4667 ( .A(n938), .Y(n4248) );
  INVX1 U4668 ( .A(n898), .Y(n4249) );
  OR2X2 U4669 ( .A(n1523), .B(n4730), .Y(n1508) );
  INVX1 U4670 ( .A(n1508), .Y(n4253) );
  INVX1 U4671 ( .A(n1508), .Y(n4254) );
  OR2X2 U4672 ( .A(n780), .B(n4381), .Y(n763) );
  INVX1 U4673 ( .A(n763), .Y(n4255) );
  INVX1 U4674 ( .A(n763), .Y(n4256) );
  INVX1 U4675 ( .A(n3749), .Y(n4257) );
  INVX1 U4676 ( .A(n3749), .Y(n4258) );
  OR2X2 U4677 ( .A(n862), .B(n4603), .Y(n851) );
  INVX1 U4678 ( .A(n851), .Y(n4259) );
  INVX1 U4679 ( .A(n851), .Y(n4260) );
  OR2X2 U4680 ( .A(n862), .B(n836), .Y(n834) );
  INVX1 U4681 ( .A(n834), .Y(n4261) );
  INVX1 U4682 ( .A(n834), .Y(n4262) );
  OR2X2 U4683 ( .A(n862), .B(n4307), .Y(n821) );
  INVX1 U4684 ( .A(n821), .Y(n4263) );
  INVX1 U4685 ( .A(n821), .Y(n4264) );
  OR2X2 U4686 ( .A(n862), .B(n4688), .Y(n804) );
  INVX1 U4687 ( .A(n804), .Y(n4265) );
  INVX1 U4688 ( .A(n804), .Y(n4266) );
  OR2X2 U4689 ( .A(n862), .B(n4308), .Y(n791) );
  INVX1 U4690 ( .A(n791), .Y(n4267) );
  INVX1 U4691 ( .A(n791), .Y(n4268) );
  OR2X2 U4692 ( .A(n862), .B(n4309), .Y(n774) );
  INVX1 U4693 ( .A(n774), .Y(n4269) );
  INVX1 U4694 ( .A(n774), .Y(n4270) );
  OR2X2 U4695 ( .A(n862), .B(n4310), .Y(n759) );
  INVX1 U4696 ( .A(n759), .Y(n4271) );
  INVX1 U4697 ( .A(n759), .Y(n4272) );
  OR2X2 U4698 ( .A(n502), .B(n4401), .Y(n456) );
  INVX1 U4699 ( .A(n456), .Y(n4273) );
  INVX1 U4700 ( .A(n2978), .Y(n4274) );
  INVX1 U4701 ( .A(n4274), .Y(n4275) );
  OR2X2 U4702 ( .A(n1665), .B(n4668), .Y(n1654) );
  INVX1 U4703 ( .A(n1654), .Y(n4276) );
  INVX1 U4704 ( .A(n1647), .Y(n4277) );
  BUFX2 U4705 ( .A(n2926), .Y(n4278) );
  INVX1 U4706 ( .A(n1382), .Y(n4279) );
  INVX1 U4707 ( .A(n1382), .Y(n4280) );
  OR2X2 U4708 ( .A(n4317), .B(n1274), .Y(n1272) );
  INVX1 U4709 ( .A(n1272), .Y(n4281) );
  INVX1 U4710 ( .A(n1072), .Y(n4282) );
  INVX1 U4711 ( .A(n1024), .Y(n4283) );
  INVX1 U4712 ( .A(n1024), .Y(n4284) );
  INVX1 U4713 ( .A(n750), .Y(n4285) );
  INVX1 U4714 ( .A(n750), .Y(n4286) );
  OR2X2 U4715 ( .A(n324), .B(n4628), .Y(n280) );
  INVX1 U4716 ( .A(n280), .Y(n4287) );
  OR2X2 U4717 ( .A(n3393), .B(n324), .Y(n258) );
  INVX1 U4718 ( .A(n258), .Y(n4288) );
  BUFX2 U4719 ( .A(n3504), .Y(n4289) );
  BUFX2 U4720 ( .A(n3506), .Y(n4290) );
  INVX1 U4721 ( .A(n1840), .Y(n4291) );
  AND2X2 U4722 ( .A(n4168), .B(n3722), .Y(n1897) );
  INVX1 U4723 ( .A(n1897), .Y(n4292) );
  AND2X2 U4724 ( .A(n4148), .B(n1886), .Y(n1875) );
  INVX1 U4725 ( .A(n1875), .Y(n4293) );
  AND2X2 U4726 ( .A(n4701), .B(n1886), .Y(n1862) );
  INVX1 U4727 ( .A(n1862), .Y(n4294) );
  AND2X2 U4728 ( .A(n1886), .B(n3262), .Y(n1851) );
  INVX1 U4729 ( .A(n1851), .Y(n4295) );
  AND2X2 U4730 ( .A(n3248), .B(n1727), .Y(n1705) );
  INVX1 U4731 ( .A(n1705), .Y(n4296) );
  AND2X2 U4732 ( .A(n2229), .B(n3724), .Y(n1560) );
  INVX1 U4733 ( .A(n1560), .Y(n4297) );
  AND2X2 U4734 ( .A(n2227), .B(n1547), .Y(n1534) );
  INVX1 U4735 ( .A(n1534), .Y(n4298) );
  AND2X2 U4736 ( .A(n4710), .B(n1547), .Y(n1519) );
  INVX1 U4737 ( .A(n1519), .Y(n4299) );
  INVX1 U4738 ( .A(n1506), .Y(n4300) );
  AND2X2 U4739 ( .A(n1547), .B(n4253), .Y(n1506) );
  AND2X2 U4740 ( .A(n3292), .B(n1208), .Y(n1184) );
  INVX1 U4741 ( .A(n1184), .Y(n4301) );
  AND2X2 U4742 ( .A(n2189), .B(n3283), .Y(n1127) );
  INVX1 U4743 ( .A(n1127), .Y(n4302) );
  AND2X2 U4744 ( .A(n2187), .B(n1112), .Y(n1101) );
  INVX1 U4745 ( .A(n1101), .Y(n4303) );
  AND2X2 U4746 ( .A(n3284), .B(n4181), .Y(n1079) );
  INVX1 U4747 ( .A(n1079), .Y(n4304) );
  AND2X2 U4748 ( .A(n3752), .B(n3052), .Y(n1053) );
  INVX1 U4749 ( .A(n1053), .Y(n4305) );
  AND2X2 U4750 ( .A(n4536), .B(n1020), .Y(n994) );
  INVX1 U4751 ( .A(n994), .Y(n4306) );
  AND2X2 U4752 ( .A(n3286), .B(n827), .Y(n823) );
  INVX1 U4753 ( .A(n823), .Y(n4307) );
  AND2X2 U4754 ( .A(n795), .B(n808), .Y(n793) );
  INVX1 U4755 ( .A(n793), .Y(n4308) );
  AND2X2 U4756 ( .A(n4595), .B(n808), .Y(n776) );
  INVX1 U4757 ( .A(n776), .Y(n4309) );
  AND2X2 U4758 ( .A(n808), .B(n4255), .Y(n761) );
  INVX1 U4759 ( .A(n761), .Y(n4310) );
  INVX1 U4760 ( .A(n506), .Y(n4311) );
  AND2X2 U4761 ( .A(n4545), .B(n4705), .Y(n436) );
  INVX1 U4762 ( .A(n436), .Y(n4312) );
  AND2X2 U4763 ( .A(n4783), .B(n3287), .Y(n207) );
  INVX1 U4764 ( .A(n207), .Y(n4313) );
  INVX1 U4765 ( .A(n1825), .Y(n4314) );
  INVX1 U4766 ( .A(n1765), .Y(n4315) );
  INVX1 U4767 ( .A(n1294), .Y(n4317) );
  INVX1 U4768 ( .A(n1294), .Y(n4318) );
  INVX1 U4769 ( .A(n918), .Y(n4319) );
  INVX1 U4770 ( .A(n708), .Y(n4320) );
  INVX1 U4771 ( .A(n1902), .Y(n4322) );
  BUFX2 U4772 ( .A(n3467), .Y(n4323) );
  AND2X2 U4773 ( .A(n3110), .B(n4589), .Y(n584) );
  INVX1 U4774 ( .A(n584), .Y(n4324) );
  INVX1 U4775 ( .A(n1719), .Y(n4325) );
  INVX1 U4776 ( .A(n2082), .Y(n4326) );
  INVX1 U4777 ( .A(n3025), .Y(n4327) );
  INVX1 U4778 ( .A(n4327), .Y(n4328) );
  INVX1 U4779 ( .A(n728), .Y(n4329) );
  BUFX2 U4780 ( .A(n3268), .Y(n4330) );
  INVX1 U4781 ( .A(n1885), .Y(n4332) );
  INVX1 U4782 ( .A(n4332), .Y(n4333) );
  INVX1 U4783 ( .A(n4332), .Y(n4334) );
  INVX1 U4784 ( .A(n1728), .Y(n4335) );
  INVX1 U4785 ( .A(n1548), .Y(n4336) );
  INVX1 U4786 ( .A(n1209), .Y(n4337) );
  INVX1 U4787 ( .A(n1021), .Y(n4338) );
  INVX1 U4788 ( .A(n807), .Y(n4339) );
  INVX1 U4789 ( .A(n4339), .Y(n4340) );
  INVX1 U4790 ( .A(n4339), .Y(n4341) );
  INVX1 U4791 ( .A(n461), .Y(n4342) );
  INVX1 U4792 ( .A(n285), .Y(n4343) );
  INVX1 U4793 ( .A(n1799), .Y(n4344) );
  AND2X2 U4794 ( .A(B[102]), .B(A[102]), .Y(n1084) );
  INVX1 U4795 ( .A(n1084), .Y(n4346) );
  INVX1 U4796 ( .A(n1084), .Y(n4347) );
  INVX1 U4797 ( .A(n1036), .Y(n4348) );
  INVX1 U4798 ( .A(n1010), .Y(n4349) );
  AND2X2 U4799 ( .A(B[110]), .B(A[110]), .Y(n986) );
  INVX1 U4800 ( .A(n986), .Y(n4350) );
  INVX1 U4801 ( .A(n986), .Y(n4351) );
  INVX1 U4802 ( .A(n828), .Y(n4352) );
  AND2X2 U4803 ( .A(B[128]), .B(A[128]), .Y(n738) );
  INVX1 U4804 ( .A(n738), .Y(n4353) );
  INVX1 U4805 ( .A(n738), .Y(n4354) );
  INVX1 U4806 ( .A(n1781), .Y(n4355) );
  INVX1 U4807 ( .A(n1699), .Y(n4356) );
  INVX1 U4808 ( .A(n2062), .Y(n4357) );
  INVX1 U4809 ( .A(n1834), .Y(n4358) );
  INVX1 U4810 ( .A(n1942), .Y(n4359) );
  INVX1 U4811 ( .A(n1635), .Y(n4360) );
  INVX1 U4812 ( .A(n1635), .Y(n4361) );
  AND2X2 U4813 ( .A(B[148]), .B(A[148]), .Y(n538) );
  INVX1 U4814 ( .A(n538), .Y(n4362) );
  INVX1 U4815 ( .A(n538), .Y(n4363) );
  INVX1 U4816 ( .A(n4367), .Y(n4364) );
  INVX1 U4817 ( .A(n4364), .Y(n4365) );
  INVX1 U4818 ( .A(n4364), .Y(n4366) );
  OR2X2 U4819 ( .A(A[156]), .B(B[156]), .Y(n4663) );
  INVX1 U4820 ( .A(n4663), .Y(n4367) );
  INVX1 U4821 ( .A(n4370), .Y(n4368) );
  INVX1 U4822 ( .A(n4368), .Y(n4369) );
  OR2X2 U4823 ( .A(A[150]), .B(B[150]), .Y(n4666) );
  INVX1 U4824 ( .A(n4666), .Y(n4370) );
  INVX1 U4825 ( .A(n4670), .Y(n4371) );
  INVX1 U4826 ( .A(n4670), .Y(n4372) );
  OR2X2 U4827 ( .A(A[146]), .B(B[146]), .Y(n4670) );
  INVX1 U4828 ( .A(n4375), .Y(n4373) );
  INVX1 U4829 ( .A(n4373), .Y(n4374) );
  OR2X2 U4830 ( .A(A[142]), .B(B[142]), .Y(n4673) );
  INVX1 U4831 ( .A(n4673), .Y(n4375) );
  INVX1 U4832 ( .A(n4379), .Y(n4376) );
  INVX1 U4833 ( .A(n4376), .Y(n4377) );
  INVX1 U4834 ( .A(n4376), .Y(n4378) );
  OR2X2 U4835 ( .A(A[116]), .B(B[116]), .Y(n4674) );
  INVX1 U4836 ( .A(n4674), .Y(n4379) );
  INVX1 U4837 ( .A(n4383), .Y(n4380) );
  INVX1 U4838 ( .A(n4380), .Y(n4381) );
  INVX1 U4839 ( .A(n4380), .Y(n4382) );
  OR2X2 U4840 ( .A(A[126]), .B(B[126]), .Y(n4675) );
  INVX1 U4841 ( .A(n4675), .Y(n4383) );
  INVX1 U4842 ( .A(n4387), .Y(n4384) );
  INVX1 U4843 ( .A(n4384), .Y(n4385) );
  INVX1 U4844 ( .A(n4384), .Y(n4386) );
  OR2X2 U4845 ( .A(A[140]), .B(B[140]), .Y(n4676) );
  INVX1 U4846 ( .A(n4676), .Y(n4387) );
  INVX1 U4847 ( .A(n4391), .Y(n4388) );
  INVX1 U4848 ( .A(n4388), .Y(n4389) );
  INVX1 U4849 ( .A(n4388), .Y(n4390) );
  OR2X2 U4850 ( .A(A[118]), .B(B[118]), .Y(n4677) );
  INVX1 U4851 ( .A(n4677), .Y(n4391) );
  INVX1 U4852 ( .A(n4394), .Y(n4392) );
  INVX1 U4853 ( .A(n4392), .Y(n4393) );
  OR2X2 U4854 ( .A(A[136]), .B(B[136]), .Y(n4697) );
  INVX1 U4855 ( .A(n4697), .Y(n4394) );
  INVX1 U4856 ( .A(n4398), .Y(n4395) );
  INVX1 U4857 ( .A(n4395), .Y(n4396) );
  INVX1 U4858 ( .A(n4395), .Y(n4397) );
  OR2X2 U4859 ( .A(A[134]), .B(B[134]), .Y(n4702) );
  INVX1 U4860 ( .A(n4702), .Y(n4398) );
  INVX1 U4861 ( .A(n4704), .Y(n4399) );
  INVX1 U4862 ( .A(n4704), .Y(n4400) );
  INVX1 U4863 ( .A(n4705), .Y(n4401) );
  INVX1 U4864 ( .A(n4405), .Y(n4402) );
  INVX1 U4865 ( .A(n4402), .Y(n4403) );
  INVX1 U4866 ( .A(n4402), .Y(n4404) );
  OR2X2 U4867 ( .A(A[14]), .B(B[14]), .Y(n4712) );
  INVX1 U4868 ( .A(n4712), .Y(n4405) );
  INVX1 U4869 ( .A(n4409), .Y(n4406) );
  INVX1 U4870 ( .A(n4406), .Y(n4407) );
  INVX1 U4871 ( .A(n4406), .Y(n4408) );
  OR2X2 U4872 ( .A(A[88]), .B(B[88]), .Y(n4713) );
  INVX1 U4873 ( .A(n4713), .Y(n4409) );
  INVX1 U4874 ( .A(n4413), .Y(n4410) );
  INVX1 U4875 ( .A(n4410), .Y(n4411) );
  INVX1 U4876 ( .A(n4410), .Y(n4412) );
  OR2X2 U4877 ( .A(A[84]), .B(B[84]), .Y(n4715) );
  INVX1 U4878 ( .A(n4715), .Y(n4413) );
  INVX1 U4879 ( .A(n4417), .Y(n4414) );
  INVX1 U4880 ( .A(n4414), .Y(n4415) );
  INVX1 U4881 ( .A(n4414), .Y(n4416) );
  OR2X2 U4882 ( .A(A[138]), .B(B[138]), .Y(n4720) );
  INVX1 U4883 ( .A(n4720), .Y(n4417) );
  INVX1 U4884 ( .A(n4421), .Y(n4418) );
  INVX1 U4885 ( .A(n4418), .Y(n4419) );
  INVX1 U4886 ( .A(n4418), .Y(n4420) );
  OR2X2 U4887 ( .A(A[130]), .B(B[130]), .Y(n4724) );
  INVX1 U4888 ( .A(n4724), .Y(n4421) );
  INVX1 U4889 ( .A(n4425), .Y(n4422) );
  INVX1 U4890 ( .A(n4422), .Y(n4423) );
  INVX1 U4891 ( .A(n4422), .Y(n4424) );
  OR2X2 U4892 ( .A(A[30]), .B(B[30]), .Y(n4732) );
  INVX1 U4893 ( .A(n4732), .Y(n4425) );
  INVX1 U4894 ( .A(n4429), .Y(n4426) );
  INVX1 U4895 ( .A(n4426), .Y(n4427) );
  INVX1 U4896 ( .A(n4426), .Y(n4428) );
  OR2X2 U4897 ( .A(A[86]), .B(B[86]), .Y(n4736) );
  INVX1 U4898 ( .A(n4736), .Y(n4429) );
  INVX1 U4899 ( .A(n4737), .Y(n4430) );
  INVX1 U4900 ( .A(n4737), .Y(n4431) );
  OR2X2 U4901 ( .A(A[80]), .B(B[80]), .Y(n4737) );
  INVX1 U4902 ( .A(n4747), .Y(n4432) );
  INVX1 U4903 ( .A(n4747), .Y(n4433) );
  OR2X2 U4904 ( .A(A[82]), .B(B[82]), .Y(n4747) );
  INVX1 U4905 ( .A(n4758), .Y(n4434) );
  INVX1 U4906 ( .A(n4758), .Y(n4435) );
  INVX1 U4907 ( .A(n4439), .Y(n4436) );
  INVX1 U4908 ( .A(n4436), .Y(n4437) );
  INVX1 U4909 ( .A(n4436), .Y(n4438) );
  OR2X2 U4910 ( .A(A[92]), .B(B[92]), .Y(n4760) );
  INVX1 U4911 ( .A(n4760), .Y(n4439) );
  INVX1 U4912 ( .A(n4443), .Y(n4440) );
  INVX1 U4913 ( .A(n4440), .Y(n4441) );
  INVX1 U4914 ( .A(n4440), .Y(n4442) );
  OR2X2 U4915 ( .A(A[70]), .B(B[70]), .Y(n4761) );
  INVX1 U4916 ( .A(n4761), .Y(n4443) );
  INVX1 U4917 ( .A(n4447), .Y(n4444) );
  INVX1 U4918 ( .A(n4444), .Y(n4445) );
  INVX1 U4919 ( .A(n4444), .Y(n4446) );
  OR2X2 U4920 ( .A(A[68]), .B(B[68]), .Y(n4762) );
  INVX1 U4921 ( .A(n4762), .Y(n4447) );
  INVX1 U4922 ( .A(n2964), .Y(n4448) );
  INVX1 U4923 ( .A(n1649), .Y(n4449) );
  INVX1 U4924 ( .A(n1649), .Y(n4450) );
  INVX1 U4925 ( .A(n2232), .Y(n4451) );
  INVX1 U4926 ( .A(n1579), .Y(n4452) );
  INVX1 U4927 ( .A(n1499), .Y(n4453) );
  INVX1 U4928 ( .A(n1499), .Y(n4454) );
  INVX1 U4929 ( .A(n4174), .Y(n4455) );
  INVX1 U4930 ( .A(n1426), .Y(n4456) );
  INVX1 U4931 ( .A(n1426), .Y(n4457) );
  INVX1 U4932 ( .A(n1384), .Y(n4459) );
  INVX1 U4933 ( .A(n4178), .Y(n4460) );
  INVX1 U4934 ( .A(n926), .Y(n4461) );
  INVX1 U4935 ( .A(n4185), .Y(n4462) );
  INVX1 U4936 ( .A(n752), .Y(n4463) );
  INVX1 U4937 ( .A(n3097), .Y(n4464) );
  INVX1 U4938 ( .A(n4464), .Y(n4465) );
  INVX1 U4939 ( .A(n654), .Y(n4466) );
  INVX1 U4940 ( .A(n614), .Y(n4467) );
  INVX1 U4941 ( .A(n4471), .Y(n4468) );
  INVX1 U4942 ( .A(n4468), .Y(n4469) );
  INVX1 U4943 ( .A(n4468), .Y(n4470) );
  OR2X2 U4944 ( .A(A[132]), .B(B[132]), .Y(n4706) );
  INVX1 U4945 ( .A(n4706), .Y(n4471) );
  INVX1 U4946 ( .A(n2268), .Y(n4472) );
  INVX1 U4947 ( .A(n2971), .Y(n4473) );
  INVX1 U4948 ( .A(n4473), .Y(n4474) );
  INVX1 U4949 ( .A(n1870), .Y(n4475) );
  INVX1 U4950 ( .A(n1791), .Y(n4476) );
  INVX1 U4951 ( .A(n1733), .Y(n4478) );
  INVX1 U4952 ( .A(n2240), .Y(n4479) );
  INVX1 U4953 ( .A(n1553), .Y(n4481) );
  INVX1 U4954 ( .A(n1553), .Y(n4482) );
  INVX1 U4955 ( .A(n2226), .Y(n4483) );
  INVX1 U4956 ( .A(n1444), .Y(n4484) );
  INVX1 U4957 ( .A(n1444), .Y(n4485) );
  INVX1 U4958 ( .A(n1320), .Y(n4486) );
  INVX1 U4959 ( .A(n1320), .Y(n4487) );
  OR2X2 U4960 ( .A(A[85]), .B(B[85]), .Y(n1278) );
  INVX1 U4961 ( .A(n1278), .Y(n4488) );
  INVX1 U4962 ( .A(n1278), .Y(n4489) );
  INVX1 U4963 ( .A(n1234), .Y(n4490) );
  INVX1 U4964 ( .A(n4247), .Y(n4491) );
  INVX1 U4965 ( .A(n1122), .Y(n4492) );
  INVX1 U4966 ( .A(n4180), .Y(n4493) );
  INVX1 U4967 ( .A(n1048), .Y(n4494) );
  INVX1 U4968 ( .A(n1048), .Y(n4495) );
  INVX1 U4969 ( .A(n2180), .Y(n4496) );
  INVX1 U4970 ( .A(n898), .Y(n4498) );
  INVX1 U4971 ( .A(n844), .Y(n4499) );
  INVX1 U4972 ( .A(n844), .Y(n4500) );
  INVX1 U4973 ( .A(n814), .Y(n4501) );
  INVX1 U4974 ( .A(n814), .Y(n4502) );
  INVX1 U4975 ( .A(n784), .Y(n4503) );
  INVX1 U4976 ( .A(n732), .Y(n4504) );
  INVX1 U4977 ( .A(n732), .Y(n4505) );
  INVX1 U4978 ( .A(n4250), .Y(n4506) );
  INVX1 U4979 ( .A(n572), .Y(n4507) );
  OR2X2 U4980 ( .A(A[147]), .B(B[147]), .Y(n554) );
  INVX1 U4981 ( .A(n554), .Y(n4508) );
  INVX1 U4982 ( .A(n554), .Y(n4509) );
  INVX1 U4983 ( .A(n530), .Y(n4510) );
  INVX1 U4984 ( .A(n530), .Y(n4511) );
  OR2X2 U4985 ( .A(A[151]), .B(B[151]), .Y(n510) );
  INVX1 U4986 ( .A(n510), .Y(n4512) );
  INVX1 U4987 ( .A(n510), .Y(n4513) );
  INVX1 U4988 ( .A(n3115), .Y(n4514) );
  INVX1 U4989 ( .A(n4514), .Y(n4515) );
  INVX1 U4990 ( .A(n466), .Y(n4516) );
  INVX1 U4991 ( .A(n466), .Y(n4517) );
  INVX1 U4992 ( .A(n420), .Y(n4518) );
  INVX1 U4993 ( .A(n420), .Y(n4519) );
  INVX1 U4994 ( .A(n396), .Y(n4520) );
  INVX1 U4995 ( .A(n396), .Y(n4521) );
  INVX1 U4996 ( .A(n378), .Y(n4522) );
  INVX1 U4997 ( .A(n354), .Y(n4523) );
  INVX1 U4998 ( .A(n3132), .Y(n4524) );
  INVX1 U4999 ( .A(n4524), .Y(n4525) );
  INVX1 U5000 ( .A(n310), .Y(n4526) );
  INVX1 U5001 ( .A(n310), .Y(n4527) );
  INVX1 U5002 ( .A(n290), .Y(n4528) );
  INVX1 U5003 ( .A(n244), .Y(n4529) );
  INVX1 U5004 ( .A(n220), .Y(n4530) );
  INVX1 U5005 ( .A(n1621), .Y(n4531) );
  INVX1 U5006 ( .A(n1621), .Y(n4532) );
  INVX1 U5007 ( .A(n1398), .Y(n4533) );
  INVX1 U5008 ( .A(n1398), .Y(n4534) );
  INVX1 U5009 ( .A(n3064), .Y(n4535) );
  INVX1 U5010 ( .A(n4535), .Y(n4536) );
  INVX1 U5011 ( .A(n3077), .Y(n4537) );
  INVX1 U5012 ( .A(n4537), .Y(n4538) );
  INVX1 U5013 ( .A(n692), .Y(n4539) );
  INVX1 U5014 ( .A(n692), .Y(n4540) );
  INVX1 U5015 ( .A(n650), .Y(n4541) );
  INVX1 U5016 ( .A(n650), .Y(n4542) );
  INVX1 U5017 ( .A(n610), .Y(n4543) );
  INVX1 U5018 ( .A(n568), .Y(n4544) );
  INVX1 U5019 ( .A(n438), .Y(n4545) );
  INVX1 U5020 ( .A(n3124), .Y(n4546) );
  INVX1 U5021 ( .A(n4546), .Y(n4547) );
  INVX1 U5022 ( .A(n3138), .Y(n4548) );
  INVX1 U5023 ( .A(n4548), .Y(n4549) );
  BUFX2 U5024 ( .A(n2915), .Y(n4550) );
  BUFX2 U5025 ( .A(n3469), .Y(n4551) );
  INVX1 U5026 ( .A(n1513), .Y(n4552) );
  BUFX2 U5027 ( .A(n2922), .Y(n4553) );
  BUFX2 U5028 ( .A(n3515), .Y(n4554) );
  INVX1 U5029 ( .A(n3751), .Y(n4555) );
  INVX1 U5030 ( .A(n3751), .Y(n4556) );
  BUFX2 U5031 ( .A(n3477), .Y(n4557) );
  INVX1 U5032 ( .A(n938), .Y(n4558) );
  BUFX2 U5033 ( .A(n3517), .Y(n4559) );
  BUFX2 U5034 ( .A(n3481), .Y(n4560) );
  BUFX2 U5035 ( .A(n3519), .Y(n4561) );
  BUFX2 U5036 ( .A(n3521), .Y(n4562) );
  BUFX2 U5037 ( .A(n3483), .Y(n4563) );
  AND2X2 U5038 ( .A(B[144]), .B(A[144]), .Y(n580) );
  INVX1 U5039 ( .A(n580), .Y(n4564) );
  INVX1 U5040 ( .A(n580), .Y(n4565) );
  AND2X2 U5041 ( .A(B[152]), .B(A[152]), .Y(n494) );
  INVX1 U5042 ( .A(n494), .Y(n4566) );
  INVX1 U5043 ( .A(n494), .Y(n4567) );
  AND2X2 U5044 ( .A(B[154]), .B(A[154]), .Y(n474) );
  INVX1 U5045 ( .A(n474), .Y(n4568) );
  INVX1 U5046 ( .A(n474), .Y(n4569) );
  INVX1 U5047 ( .A(n450), .Y(n4570) );
  INVX1 U5048 ( .A(n450), .Y(n4571) );
  AND2X2 U5049 ( .A(B[158]), .B(A[158]), .Y(n428) );
  INVX1 U5050 ( .A(n428), .Y(n4572) );
  INVX1 U5051 ( .A(n428), .Y(n4573) );
  AND2X2 U5052 ( .A(B[160]), .B(A[160]), .Y(n404) );
  INVX1 U5053 ( .A(n404), .Y(n4574) );
  INVX1 U5054 ( .A(n404), .Y(n4575) );
  INVX1 U5055 ( .A(n298), .Y(n4576) );
  INVX1 U5056 ( .A(n252), .Y(n4577) );
  INVX1 U5057 ( .A(n1018), .Y(n4578) );
  INVX1 U5058 ( .A(n1018), .Y(n4579) );
  INVX1 U5059 ( .A(n3528), .Y(n4580) );
  INVX1 U5060 ( .A(n4580), .Y(n4581) );
  INVX1 U5061 ( .A(n921), .Y(n4582) );
  INVX1 U5062 ( .A(n711), .Y(n4583) );
  INVX1 U5063 ( .A(n4682), .Y(n4584) );
  INVX1 U5064 ( .A(n545), .Y(n4585) );
  INVX1 U5065 ( .A(n369), .Y(n4586) );
  INVX1 U5066 ( .A(n3103), .Y(n4587) );
  INVX1 U5067 ( .A(n4587), .Y(n4588) );
  INVX1 U5068 ( .A(n668), .Y(n4589) );
  INVX1 U5069 ( .A(n668), .Y(n4590) );
  INVX1 U5070 ( .A(n1663), .Y(n4591) );
  INVX1 U5071 ( .A(n1663), .Y(n4592) );
  INVX1 U5072 ( .A(n778), .Y(n4593) );
  INVX1 U5073 ( .A(n778), .Y(n4594) );
  INVX1 U5074 ( .A(n778), .Y(n4595) );
  INVX1 U5075 ( .A(n500), .Y(n4596) );
  INVX1 U5076 ( .A(n500), .Y(n4597) );
  INVX1 U5077 ( .A(n324), .Y(n4598) );
  INVX1 U5078 ( .A(n324), .Y(n4599) );
  INVX1 U5079 ( .A(n1149), .Y(n4600) );
  INVX1 U5080 ( .A(n1149), .Y(n4601) );
  INVX1 U5081 ( .A(n853), .Y(n4602) );
  INVX1 U5082 ( .A(n853), .Y(n4603) );
  INVX1 U5083 ( .A(n577), .Y(n4604) );
  INVX1 U5084 ( .A(n577), .Y(n4605) );
  INVX1 U5085 ( .A(n535), .Y(n4606) );
  INVX1 U5086 ( .A(n535), .Y(n4607) );
  INVX1 U5087 ( .A(n535), .Y(n4608) );
  INVX1 U5088 ( .A(n491), .Y(n4609) );
  INVX1 U5089 ( .A(n491), .Y(n4610) );
  INVX1 U5090 ( .A(n471), .Y(n4611) );
  INVX1 U5091 ( .A(n471), .Y(n4612) );
  INVX1 U5092 ( .A(n425), .Y(n4613) );
  INVX1 U5093 ( .A(n425), .Y(n4614) );
  INVX1 U5094 ( .A(n401), .Y(n4615) );
  INVX1 U5095 ( .A(n401), .Y(n4616) );
  INVX1 U5096 ( .A(n383), .Y(n4617) );
  INVX1 U5097 ( .A(n383), .Y(n4618) );
  INVX1 U5098 ( .A(n359), .Y(n4619) );
  INVX1 U5099 ( .A(n339), .Y(n4620) );
  INVX1 U5100 ( .A(n339), .Y(n4621) );
  INVX1 U5101 ( .A(n339), .Y(n4622) );
  INVX1 U5102 ( .A(n315), .Y(n4623) );
  INVX1 U5103 ( .A(n315), .Y(n4624) );
  INVX1 U5104 ( .A(n295), .Y(n4625) );
  INVX1 U5105 ( .A(n295), .Y(n4626) );
  INVX1 U5106 ( .A(n282), .Y(n4627) );
  INVX1 U5107 ( .A(n282), .Y(n4628) );
  INVX1 U5108 ( .A(n271), .Y(n4629) );
  INVX1 U5109 ( .A(n271), .Y(n4630) );
  INVX1 U5110 ( .A(n249), .Y(n4631) );
  INVX1 U5111 ( .A(n249), .Y(n4632) );
  INVX1 U5112 ( .A(n225), .Y(n4633) );
  INVX1 U5113 ( .A(n1926), .Y(n4635) );
  INVX1 U5114 ( .A(n862), .Y(n4636) );
  INVX4 U5115 ( .A(n15), .Y(n4652) );
  XNOR2X1 U5116 ( .A(n3583), .B(n4638), .Y(SUM[155]) );
  AND2X2 U5117 ( .A(n4165), .B(n2132), .Y(n4638) );
  INVX1 U5118 ( .A(n4746), .Y(n4639) );
  BUFX2 U5119 ( .A(n3726), .Y(n4640) );
  INVX1 U5120 ( .A(n2843), .Y(n4641) );
  INVX1 U5121 ( .A(n4641), .Y(n4642) );
  XNOR2X1 U5122 ( .A(n3577), .B(n4644), .Y(SUM[26]) );
  AND2X2 U5123 ( .A(n4322), .B(n4168), .Y(n4644) );
  XOR2X1 U5124 ( .A(n1720), .B(n4645), .Y(SUM[44]) );
  AND2X2 U5125 ( .A(n2997), .B(n4170), .Y(n4645) );
  INVX1 U5126 ( .A(n1819), .Y(n4646) );
  XNOR2X1 U5127 ( .A(n3500), .B(n4647), .Y(SUM[4]) );
  AND2X2 U5128 ( .A(n3893), .B(n2091), .Y(n4647) );
  XNOR2X1 U5129 ( .A(n196), .B(n4777), .Y(SUM[1]) );
  XNOR2X1 U5130 ( .A(n3578), .B(n4648), .Y(SUM[27]) );
  AND2X2 U5131 ( .A(n2977), .B(n2260), .Y(n4648) );
  XNOR2X1 U5132 ( .A(n2064), .B(n4649), .Y(SUM[8]) );
  AND2X2 U5133 ( .A(n3497), .B(n2062), .Y(n4649) );
  INVX1 U5134 ( .A(n3527), .Y(n4650) );
  INVX1 U5135 ( .A(n4650), .Y(n4651) );
  XNOR2X1 U5136 ( .A(n3580), .B(n4653), .Y(SUM[142]) );
  AND2X2 U5137 ( .A(n3487), .B(n4373), .Y(n4653) );
  XNOR2X1 U5138 ( .A(n3581), .B(n4654), .Y(SUM[148]) );
  AND2X2 U5139 ( .A(n4363), .B(n2139), .Y(n4654) );
  XNOR2X1 U5140 ( .A(n3582), .B(n4655), .Y(SUM[150]) );
  AND2X2 U5141 ( .A(n3112), .B(n2137), .Y(n4655) );
  XNOR2X1 U5142 ( .A(n3585), .B(n4656), .Y(SUM[166]) );
  AND2X2 U5143 ( .A(n2918), .B(n2121), .Y(n4656) );
  XNOR2X1 U5144 ( .A(n3584), .B(n4657), .Y(SUM[163]) );
  AND2X2 U5145 ( .A(n3126), .B(n378), .Y(n4657) );
  XNOR2X1 U5146 ( .A(n3586), .B(n4658), .Y(SUM[168]) );
  AND2X2 U5147 ( .A(n3491), .B(n2119), .Y(n4658) );
  INVX1 U5148 ( .A(n4773), .Y(n4659) );
  INVX1 U5149 ( .A(n944), .Y(n4660) );
  INVX1 U5150 ( .A(n1919), .Y(n4661) );
  BUFX2 U5151 ( .A(n3465), .Y(n4662) );
  INVX1 U5152 ( .A(n4771), .Y(n4664) );
  INVX1 U5153 ( .A(n1424), .Y(n4665) );
  INVX4 U5154 ( .A(n4773), .Y(n4774) );
  INVX1 U5155 ( .A(n1927), .Y(n4667) );
  INVX1 U5156 ( .A(n1656), .Y(n4668) );
  INVX1 U5157 ( .A(n1251), .Y(n4669) );
  INVX1 U5158 ( .A(n729), .Y(n4672) );
  AND2X2 U5159 ( .A(B[10]), .B(A[10]), .Y(n4678) );
  INVX1 U5160 ( .A(n4754), .Y(n4679) );
  BUFX2 U5161 ( .A(n3501), .Y(n4680) );
  INVX1 U5162 ( .A(n587), .Y(n4681) );
  INVX1 U5163 ( .A(n4681), .Y(n4682) );
  INVX1 U5164 ( .A(n4681), .Y(n4683) );
  INVX1 U5165 ( .A(n4681), .Y(n4684) );
  INVX1 U5166 ( .A(n2074), .Y(n4686) );
  INVX2 U5167 ( .A(n4685), .Y(n2072) );
  OAI21X1 U5168 ( .A(n3500), .B(n4687), .C(n4686), .Y(n4685) );
  OR2X2 U5169 ( .A(n2082), .B(n2075), .Y(n4687) );
  INVX1 U5170 ( .A(n808), .Y(n4688) );
  AND2X2 U5171 ( .A(n3729), .B(n2841), .Y(n4689) );
  INVX8 U5172 ( .A(n4698), .Y(n4794) );
  INVX1 U5173 ( .A(n2868), .Y(n4690) );
  INVX1 U5174 ( .A(n4690), .Y(n4691) );
  OR2X2 U5175 ( .A(A[7]), .B(B[7]), .Y(n4692) );
  INVX1 U5176 ( .A(n1493), .Y(n4693) );
  OR2X2 U5177 ( .A(A[6]), .B(B[6]), .Y(n4694) );
  INVX1 U5178 ( .A(n4694), .Y(n2075) );
  INVX4 U5179 ( .A(n2910), .Y(n4776) );
  INVX4 U5180 ( .A(n2909), .Y(n4775) );
  XOR2X1 U5181 ( .A(n1636), .B(n4696), .Y(SUM[52]) );
  AND2X2 U5182 ( .A(n4361), .B(n1632), .Y(n4696) );
  BUFX2 U5183 ( .A(n3505), .Y(n4786) );
  AND2X2 U5184 ( .A(n2895), .B(n3283), .Y(n1134) );
  BUFX2 U5185 ( .A(n3725), .Y(n4699) );
  INVX1 U5186 ( .A(n1970), .Y(n4700) );
  INVX1 U5187 ( .A(n1866), .Y(n4701) );
  INVX1 U5188 ( .A(n1632), .Y(n4703) );
  INVX1 U5189 ( .A(n1476), .Y(n4707) );
  AND2X2 U5190 ( .A(n3244), .B(n3265), .Y(n4708) );
  INVX1 U5191 ( .A(n4708), .Y(n1340) );
  INVX1 U5192 ( .A(n1682), .Y(n4709) );
  INVX1 U5193 ( .A(n1523), .Y(n4710) );
  INVX1 U5194 ( .A(n2231), .Y(n4711) );
  AND2X2 U5195 ( .A(n3249), .B(n3278), .Y(n4714) );
  INVX1 U5196 ( .A(n4714), .Y(n1456) );
  INVX1 U5197 ( .A(n4708), .Y(n4716) );
  INVX1 U5198 ( .A(n967), .Y(n4717) );
  INVX1 U5199 ( .A(n4717), .Y(n4718) );
  INVX1 U5200 ( .A(n4717), .Y(n4719) );
  OR2X2 U5201 ( .A(A[0]), .B(B[0]), .Y(n4784) );
  INVX4 U5202 ( .A(n4786), .Y(n1335) );
  INVX1 U5203 ( .A(n4173), .Y(n4721) );
  INVX1 U5204 ( .A(n4719), .Y(n4722) );
  INVX1 U5205 ( .A(n3739), .Y(n967) );
  INVX1 U5206 ( .A(n1112), .Y(n4723) );
  XNOR2X1 U5207 ( .A(n2072), .B(n4725), .Y(SUM[7]) );
  AND2X2 U5208 ( .A(n2960), .B(n4692), .Y(n4725) );
  INVX1 U5209 ( .A(n1967), .Y(n4726) );
  INVX1 U5210 ( .A(n1219), .Y(n4729) );
  BUFX4 U5211 ( .A(n1155), .Y(n4787) );
  INVX1 U5212 ( .A(n2225), .Y(n4730) );
  INVX1 U5213 ( .A(n1596), .Y(n4731) );
  INVX1 U5214 ( .A(n4146), .Y(n4733) );
  INVX1 U5215 ( .A(n4759), .Y(n4734) );
  XOR2X1 U5216 ( .A(n2050), .B(n4735), .Y(SUM[10]) );
  AND2X2 U5217 ( .A(n3509), .B(n2048), .Y(n4735) );
  INVX1 U5218 ( .A(n1595), .Y(n4739) );
  BUFX2 U5219 ( .A(n2839), .Y(n4740) );
  BUFX2 U5220 ( .A(n407), .Y(n4741) );
  INVX1 U5221 ( .A(n1547), .Y(n4742) );
  OR2X2 U5222 ( .A(A[1]), .B(B[1]), .Y(n4743) );
  OR2X2 U5223 ( .A(n4324), .B(n3123), .Y(n4781) );
  INVX4 U5224 ( .A(n4781), .Y(n406) );
  INVX1 U5225 ( .A(n671), .Y(n4744) );
  XNOR2X1 U5226 ( .A(n3575), .B(n4745), .Y(SUM[5]) );
  AND2X2 U5227 ( .A(n2958), .B(n2282), .Y(n4745) );
  OR2X2 U5228 ( .A(A[2]), .B(B[2]), .Y(n4746) );
  XNOR2X1 U5229 ( .A(n4749), .B(n4748), .Y(SUM[18]) );
  OAI21X1 U5230 ( .A(n4728), .B(n1982), .C(n1985), .Y(n4749) );
  AND2X2 U5231 ( .A(n2966), .B(n2269), .Y(n4750) );
  INVX1 U5232 ( .A(n4144), .Y(n4751) );
  INVX1 U5233 ( .A(n1886), .Y(n4752) );
  INVX2 U5234 ( .A(n3739), .Y(n4753) );
  OR2X2 U5235 ( .A(A[9]), .B(B[9]), .Y(n4754) );
  XNOR2X1 U5236 ( .A(n3576), .B(n4755), .Y(SUM[22]) );
  AND2X2 U5237 ( .A(n2970), .B(n4146), .Y(n4755) );
  INVX1 U5238 ( .A(n4175), .Y(n4756) );
  BUFX2 U5239 ( .A(n3503), .Y(n4757) );
  OR2X2 U5240 ( .A(A[94]), .B(B[94]), .Y(n4759) );
  INVX1 U5241 ( .A(n2019), .Y(n4763) );
  INVX1 U5242 ( .A(n4792), .Y(n4764) );
  INVX1 U5243 ( .A(n2221), .Y(n4765) );
  INVX1 U5244 ( .A(n1389), .Y(n4766) );
  BUFX2 U5245 ( .A(n3502), .Y(n4767) );
  INVX1 U5246 ( .A(n1250), .Y(n4769) );
  XNOR2X1 U5247 ( .A(n3579), .B(n4770), .Y(SUM[98]) );
  AND2X2 U5248 ( .A(n4323), .B(n2189), .Y(n4770) );
  OR2X2 U5249 ( .A(A[78]), .B(B[78]), .Y(n4771) );
  INVX1 U5250 ( .A(n1208), .Y(n4772) );
  INVX1 U5251 ( .A(n7), .Y(n4773) );
  AND2X2 U5252 ( .A(n4778), .B(n4784), .Y(SUM[0]) );
  AND2X2 U5253 ( .A(n2956), .B(n4743), .Y(n196) );
  AND2X2 U5254 ( .A(B[0]), .B(A[0]), .Y(n2107) );
  INVX1 U5255 ( .A(n2852), .Y(n4777) );
  INVX1 U5256 ( .A(n2852), .Y(n4778) );
  OR2X2 U5257 ( .A(A[18]), .B(B[18]), .Y(n1977) );
  INVX1 U5258 ( .A(n1977), .Y(n4779) );
  INVX1 U5259 ( .A(n1977), .Y(n4780) );
  BUFX2 U5260 ( .A(n2839), .Y(n4790) );
  INVX1 U5261 ( .A(n3328), .Y(n230) );
  INVX1 U5262 ( .A(n3363), .Y(n234) );
  INVX1 U5263 ( .A(n3358), .Y(n320) );
  INVX1 U5264 ( .A(n3354), .Y(n344) );
  INVX1 U5265 ( .A(n2950), .Y(n254) );
  INVX1 U5266 ( .A(n3362), .Y(n276) );
  INVX1 U5267 ( .A(n3360), .Y(n300) );
  INVX1 U5268 ( .A(n3352), .Y(n364) );
  INVX1 U5269 ( .A(n3876), .Y(n1224) );
  INVX1 U5270 ( .A(n3891), .Y(n476) );
  INVX1 U5271 ( .A(n4161), .Y(n430) );
  INVX1 U5272 ( .A(n4156), .Y(n1178) );
  INVX1 U5273 ( .A(n3877), .Y(n1200) );
  INVX1 U5274 ( .A(n3378), .Y(n1244) );
  INVX1 U5275 ( .A(n3392), .Y(n520) );
  INVX1 U5276 ( .A(n3390), .Y(n540) );
  INVX1 U5277 ( .A(n3879), .Y(n496) );
  INVX1 U5278 ( .A(n3367), .Y(n1268) );
  INVX1 U5279 ( .A(n3296), .Y(n1926) );
  INVX1 U5280 ( .A(n3302), .Y(n1250) );
  INVX1 U5281 ( .A(n4597), .Y(n502) );
  INVX1 U5282 ( .A(n2906), .Y(n1765) );
  INVX1 U5283 ( .A(n4590), .Y(n670) );
  INVX1 U5284 ( .A(n3305), .Y(n1014) );
  INVX1 U5285 ( .A(n4137), .Y(n1040) );
  INVX1 U5286 ( .A(n3284), .Y(n1088) );
  INVX1 U5287 ( .A(n3306), .Y(n990) );
  INVX1 U5288 ( .A(n3272), .Y(n1783) );
  INVX1 U5289 ( .A(n993), .Y(n991) );
  INVX1 U5290 ( .A(n893), .Y(n891) );
  INVX1 U5291 ( .A(n3348), .Y(n808) );
  INVX1 U5292 ( .A(n1620), .Y(n1618) );
  INVX1 U5293 ( .A(n3734), .Y(n1643) );
  INVX1 U5294 ( .A(n4318), .Y(n1292) );
  INVX1 U5295 ( .A(n3464), .Y(n368) );
  INVX1 U5296 ( .A(n3738), .Y(n544) );
  INVX1 U5297 ( .A(n1488), .Y(n7) );
  INVX1 U5298 ( .A(n3554), .Y(n231) );
  INVX1 U5299 ( .A(n1043), .Y(n1041) );
  INVX1 U5300 ( .A(n1746), .Y(n1744) );
  INVX1 U5301 ( .A(n1091), .Y(n1089) );
  INVX1 U5302 ( .A(n1704), .Y(n1702) );
  INVX1 U5303 ( .A(n1724), .Y(n1722) );
  INVX1 U5304 ( .A(n3346), .Y(n890) );
  INVX1 U5305 ( .A(n3336), .Y(n1617) );
  INVX1 U5306 ( .A(n3350), .Y(n388) );
  INVX1 U5307 ( .A(n3374), .Y(n1354) );
  INVX1 U5308 ( .A(n3386), .Y(n606) );
  INVX1 U5309 ( .A(n4151), .Y(n1436) );
  INVX1 U5310 ( .A(n3382), .Y(n688) );
  INVX1 U5311 ( .A(n3384), .Y(n646) );
  INVX1 U5312 ( .A(n3372), .Y(n1394) );
  INVX1 U5313 ( .A(n3376), .Y(n1312) );
  INVX1 U5314 ( .A(n3388), .Y(n564) );
  INVX1 U5315 ( .A(n523), .Y(n521) );
  INVX1 U5316 ( .A(n543), .Y(n541) );
  INVX1 U5317 ( .A(n3545), .Y(n431) );
  INVX1 U5318 ( .A(n499), .Y(n497) );
  INVX1 U5319 ( .A(n567), .Y(n565) );
  INVX1 U5320 ( .A(n3544), .Y(n453) );
  INVX1 U5321 ( .A(n3542), .Y(n477) );
  INVX1 U5322 ( .A(n3538), .Y(n647) );
  INVX1 U5323 ( .A(n3530), .Y(n1395) );
  INVX1 U5324 ( .A(n1227), .Y(n1225) );
  INVX1 U5325 ( .A(n1315), .Y(n1313) );
  INVX1 U5326 ( .A(n4235), .Y(n1179) );
  INVX1 U5327 ( .A(n1247), .Y(n1245) );
  INVX1 U5328 ( .A(n1291), .Y(n1289) );
  INVX1 U5329 ( .A(n1271), .Y(n1269) );
  INVX1 U5330 ( .A(n1203), .Y(n1201) );
  INVX1 U5331 ( .A(n691), .Y(n689) );
  INVX1 U5332 ( .A(n3531), .Y(n1355) );
  INVX1 U5333 ( .A(n3539), .Y(n607) );
  INVX1 U5334 ( .A(n1439), .Y(n1437) );
  INVX1 U5335 ( .A(n1947), .Y(n1945) );
  INVX1 U5336 ( .A(n3550), .Y(n321) );
  INVX1 U5337 ( .A(n3549), .Y(n345) );
  INVX1 U5338 ( .A(n3553), .Y(n255) );
  INVX1 U5339 ( .A(n3552), .Y(n277) );
  INVX1 U5340 ( .A(n3551), .Y(n301) );
  INVX1 U5341 ( .A(n3548), .Y(n365) );
  INVX1 U5342 ( .A(n3546), .Y(n389) );
  INVX1 U5343 ( .A(n1014), .Y(n4789) );
  INVX1 U5344 ( .A(n1047), .Y(n1045) );
  INVX1 U5345 ( .A(n2858), .Y(n1748) );
  INVX1 U5346 ( .A(n1095), .Y(n1093) );
  INVX1 U5347 ( .A(n1790), .Y(n1788) );
  INVX1 U5348 ( .A(n3231), .Y(n235) );
  INVX1 U5349 ( .A(n3535), .Y(n1021) );
  INVX1 U5350 ( .A(n2857), .Y(n1728) );
  INVX1 U5351 ( .A(n4579), .Y(n1020) );
  INVX1 U5352 ( .A(n529), .Y(n527) );
  INVX1 U5353 ( .A(n3543), .Y(n461) );
  INVX1 U5354 ( .A(n485), .Y(n483) );
  INVX1 U5355 ( .A(n3541), .Y(n545) );
  INVX1 U5356 ( .A(n3533), .Y(n1209) );
  INVX1 U5357 ( .A(n1233), .Y(n1231) );
  INVX1 U5358 ( .A(n3532), .Y(n1293) );
  INVX1 U5359 ( .A(n1277), .Y(n1275) );
  INVX1 U5360 ( .A(n219), .Y(n217) );
  INVX1 U5361 ( .A(n283), .Y(n285) );
  INVX1 U5362 ( .A(n3547), .Y(n369) );
  INVX1 U5363 ( .A(n309), .Y(n307) );
  INVX1 U5364 ( .A(n353), .Y(n351) );
  INVX1 U5365 ( .A(n863), .Y(n865) );
  INVX1 U5366 ( .A(n1594), .Y(n1596) );
  INVX1 U5367 ( .A(n1574), .Y(n1572) );
  INVX1 U5368 ( .A(n1909), .Y(n1907) );
  INVX1 U5369 ( .A(n3335), .Y(n1803) );
  INVX1 U5370 ( .A(n1249), .Y(n1251) );
  INVX1 U5371 ( .A(n501), .Y(n503) );
  INVX1 U5372 ( .A(n325), .Y(n327) );
  INVX1 U5373 ( .A(n3500), .Y(n2093) );
  INVX1 U5374 ( .A(n839), .Y(n837) );
  INVX1 U5375 ( .A(n2103), .Y(n2102) );
  INVX1 U5376 ( .A(n4341), .Y(n809) );
  INVX1 U5377 ( .A(n3529), .Y(n1548) );
  INVX1 U5378 ( .A(n4334), .Y(n1887) );
  INVX1 U5379 ( .A(n4680), .Y(n2036) );
  INVX1 U5380 ( .A(n1522), .Y(n1524) );
  INVX1 U5381 ( .A(n3536), .Y(n921) );
  INVX1 U5382 ( .A(n3537), .Y(n711) );
  INVX1 U5383 ( .A(n3286), .Y(n836) );
  INVX1 U5384 ( .A(n3724), .Y(n1571) );
  INVX1 U5385 ( .A(n3283), .Y(n1136) );
  INVX1 U5386 ( .A(n3722), .Y(n1906) );
  INVX1 U5387 ( .A(n3287), .Y(n216) );
  INVX1 U5388 ( .A(n3303), .Y(n1044) );
  INVX1 U5389 ( .A(n2840), .Y(n1092) );
  INVX1 U5390 ( .A(n3281), .Y(n1230) );
  INVX1 U5391 ( .A(n3323), .Y(n482) );
  INVX1 U5392 ( .A(n3310), .Y(n526) );
  INVX1 U5393 ( .A(n3252), .Y(n1274) );
  INVX1 U5394 ( .A(n3273), .Y(n1747) );
  INVX1 U5395 ( .A(n3298), .Y(n1787) );
  INVX1 U5396 ( .A(n2988), .Y(n1823) );
  INVX1 U5397 ( .A(n3731), .Y(n2051) );
  INVX1 U5398 ( .A(n4134), .Y(n1743) );
  INVX1 U5399 ( .A(n3221), .Y(n2266) );
  INVX1 U5400 ( .A(n3404), .Y(n2260) );
  INVX1 U5401 ( .A(n4435), .Y(n2211) );
  INVX1 U5402 ( .A(n4600), .Y(n2191) );
  INVX1 U5403 ( .A(n3430), .Y(n2221) );
  INVX1 U5404 ( .A(n4780), .Y(n2269) );
  INVX1 U5405 ( .A(n3400), .Y(n2204) );
  INVX1 U5406 ( .A(n4489), .Y(n2202) );
  INVX1 U5407 ( .A(n4463), .Y(n2160) );
  INVX1 U5408 ( .A(n4499), .Y(n2166) );
  INVX1 U5409 ( .A(n3434), .Y(n2184) );
  INVX1 U5410 ( .A(n4492), .Y(n2188) );
  INVX1 U5411 ( .A(n4603), .Y(n2167) );
  INVX1 U5412 ( .A(n4400), .Y(n2173) );
  INVX1 U5413 ( .A(n3343), .Y(n2208) );
  INVX1 U5414 ( .A(n3908), .Y(n2214) );
  INVX1 U5415 ( .A(n4457), .Y(n2216) );
  INVX1 U5416 ( .A(n4474), .Y(n2264) );
  INVX1 U5417 ( .A(n2952), .Y(n2180) );
  INVX1 U5418 ( .A(n4475), .Y(n2258) );
  INVX1 U5419 ( .A(n4407), .Y(n2199) );
  INVX1 U5420 ( .A(n4432), .Y(n2205) );
  INVX1 U5421 ( .A(n4411), .Y(n2203) );
  INVX1 U5422 ( .A(n3412), .Y(n2222) );
  INVX1 U5423 ( .A(n3409), .Y(n2270) );
  INVX1 U5424 ( .A(n4430), .Y(n2207) );
  INVX1 U5425 ( .A(n3031), .Y(n2200) );
  INVX1 U5426 ( .A(n4502), .Y(n2164) );
  INVX1 U5427 ( .A(n4494), .Y(n2182) );
  INVX1 U5428 ( .A(n3345), .Y(n2176) );
  INVX1 U5429 ( .A(n4484), .Y(n2218) );
  INVX1 U5430 ( .A(n4437), .Y(n2195) );
  INVX1 U5431 ( .A(n4394), .Y(n2151) );
  INVX1 U5432 ( .A(n4605), .Y(n2143) );
  INVX1 U5433 ( .A(n4520), .Y(n2126) );
  INVX1 U5434 ( .A(n2953), .Y(n2130) );
  INVX1 U5435 ( .A(n4517), .Y(n2132) );
  INVX1 U5436 ( .A(n4519), .Y(n2128) );
  INVX1 U5437 ( .A(n4515), .Y(n2134) );
  INVX1 U5438 ( .A(n4465), .Y(n2152) );
  INVX1 U5439 ( .A(n4526), .Y(n2118) );
  INVX1 U5440 ( .A(n4525), .Y(n2120) );
  INVX1 U5441 ( .A(n4513), .Y(n2136) );
  INVX1 U5442 ( .A(n4510), .Y(n2138) );
  INVX1 U5443 ( .A(n3107), .Y(n2144) );
  INVX1 U5444 ( .A(n3101), .Y(n2148) );
  INVX1 U5445 ( .A(n3094), .Y(n2156) );
  INVX1 U5446 ( .A(n4509), .Y(n2140) );
  INVX1 U5447 ( .A(n2954), .Y(n2114) );
  INVX1 U5448 ( .A(n4633), .Y(n2111) );
  INVX1 U5449 ( .A(n3127), .Y(n2123) );
  INVX1 U5450 ( .A(n4614), .Y(n2129) );
  INVX1 U5451 ( .A(n4624), .Y(n2119) );
  INVX1 U5452 ( .A(n4621), .Y(n2121) );
  INVX1 U5453 ( .A(n4370), .Y(n2137) );
  INVX1 U5454 ( .A(n4607), .Y(n2139) );
  INVX1 U5455 ( .A(n4626), .Y(n2117) );
  INVX1 U5456 ( .A(n4610), .Y(n2135) );
  INVX1 U5457 ( .A(n4632), .Y(n2113) );
  INVX1 U5458 ( .A(n4630), .Y(n2115) );
  INVX1 U5459 ( .A(n4504), .Y(n2158) );
  INVX1 U5460 ( .A(n2968), .Y(n2268) );
  INVX1 U5461 ( .A(n3411), .Y(n2282) );
  INVX1 U5462 ( .A(n4616), .Y(n2127) );
  INVX1 U5463 ( .A(n4617), .Y(n2125) );
  INVX1 U5464 ( .A(n4611), .Y(n2133) );
  INVX1 U5465 ( .A(n4415), .Y(n2149) );
  INVX1 U5466 ( .A(n4469), .Y(n2155) );
  INVX1 U5467 ( .A(n945), .Y(n947) );
  INVX1 U5468 ( .A(n4740), .Y(n409) );
  INVX1 U5469 ( .A(n625), .Y(n627) );
  INVX1 U5470 ( .A(n1373), .Y(n1375) );
  INVX1 U5471 ( .A(n779), .Y(n781) );
  INVX1 U5472 ( .A(n4323), .Y(n1130) );
  INVX1 U5473 ( .A(n2975), .Y(n1900) );
  INVX1 U5474 ( .A(n4347), .Y(n1082) );
  INVX1 U5475 ( .A(n1865), .Y(n1867) );
  INVX1 U5476 ( .A(n4351), .Y(n984) );
  INVX1 U5477 ( .A(n1786), .Y(n1784) );
  INVX1 U5478 ( .A(n4136), .Y(n1721) );
  INVX1 U5479 ( .A(n3017), .Y(n2225) );
  INVX1 U5480 ( .A(n3396), .Y(n2231) );
  INVX1 U5481 ( .A(n4450), .Y(n2236) );
  INVX1 U5482 ( .A(n3420), .Y(n2248) );
  INVX1 U5483 ( .A(n4454), .Y(n2224) );
  INVX1 U5484 ( .A(n3406), .Y(n2242) );
  INVX1 U5485 ( .A(n3873), .Y(n1701) );
  INVX1 U5486 ( .A(n4721), .Y(n2233) );
  INVX1 U5487 ( .A(n4478), .Y(n2244) );
  INVX1 U5488 ( .A(n3422), .Y(n2240) );
  INVX1 U5489 ( .A(n4476), .Y(n2250) );
  INVX1 U5490 ( .A(n3015), .Y(n2226) );
  INVX1 U5491 ( .A(n4482), .Y(n2228) );
  INVX1 U5492 ( .A(n3005), .Y(n2232) );
  INVX1 U5493 ( .A(n4592), .Y(n1665) );
  INVX1 U5494 ( .A(n4595), .Y(n780) );
  INVX1 U5495 ( .A(n3277), .Y(n1523) );
  INVX1 U5496 ( .A(n2983), .Y(n1866) );
  INVX1 U5497 ( .A(n3270), .Y(n2019) );
  INVX1 U5498 ( .A(n406), .Y(n408) );
  INVX1 U5499 ( .A(n4330), .Y(n626) );
  INVX1 U5500 ( .A(n3279), .Y(n1476) );
  INVX1 U5501 ( .A(n3308), .Y(n728) );
  INVX1 U5502 ( .A(n3294), .Y(n2082) );
  INVX1 U5503 ( .A(n1664), .Y(n1666) );
  INVX1 U5504 ( .A(n2018), .Y(n2020) );
  INVX1 U5505 ( .A(n3555), .Y(n1819) );
  INVX1 U5506 ( .A(n2997), .Y(n1717) );
  INVX1 U5507 ( .A(n2999), .Y(n1697) );
  INVX1 U5508 ( .A(n2991), .Y(n1779) );
  INVX1 U5509 ( .A(n2990), .Y(n1797) );
  INVX1 U5510 ( .A(n3235), .Y(n795) );
  INVX1 U5511 ( .A(n3426), .Y(n2227) );
  INVX1 U5512 ( .A(n3233), .Y(n2187) );
  INVX1 U5513 ( .A(n3043), .Y(n2189) );
  INVX1 U5514 ( .A(n3338), .Y(n2229) );
  INVX1 U5515 ( .A(n3419), .Y(n2251) );
  INVX1 U5516 ( .A(n3369), .Y(n2253) );
  INVX1 U5517 ( .A(n4142), .Y(n210) );
  INVX1 U5518 ( .A(n204), .Y(n202) );
  INVX1 U5519 ( .A(n4354), .Y(n736) );
  INVX1 U5520 ( .A(n3414), .Y(n2275) );
  OR2X1 U5521 ( .A(A[178]), .B(B[178]), .Y(n4783) );
  OR2X1 U5522 ( .A(A[179]), .B(B[179]), .Y(n4785) );
  INVX1 U5523 ( .A(n3534), .Y(n1113) );
  INVX1 U5524 ( .A(n727), .Y(n729) );
  INVX1 U5525 ( .A(n3334), .Y(n1886) );
  INVX1 U5526 ( .A(n3340), .Y(n1547) );
  INVX1 U5527 ( .A(n1139), .Y(n1137) );
  INVX1 U5528 ( .A(n2893), .Y(n1067) );
  INVX1 U5529 ( .A(n3736), .Y(n1112) );
  INVX1 U5530 ( .A(n3540), .Y(n587) );
  INVX1 U5531 ( .A(n3331), .Y(n2035) );
  INVX1 U5532 ( .A(n669), .Y(n671) );
  INVX1 U5533 ( .A(n2054), .Y(n2052) );
  INVX1 U5534 ( .A(n2081), .Y(n2083) );
  INVX1 U5535 ( .A(n3525), .Y(n1967) );
  INVX1 U5536 ( .A(n3431), .Y(n1208) );
  INVX1 U5537 ( .A(n1983), .Y(n1985) );
  INVX1 U5538 ( .A(n1925), .Y(n1927) );
  INVX1 U5539 ( .A(n4767), .Y(n1804) );
  INVX1 U5540 ( .A(n3725), .Y(n1727) );
  INVX1 U5541 ( .A(n4788), .Y(n1013) );
  AOI21X1 U5542 ( .A(n4789), .B(n2875), .C(n1017), .Y(n4788) );
  INVX1 U5543 ( .A(n2897), .Y(n1824) );
  INVX1 U5544 ( .A(n3473), .Y(n1484) );
  INVX1 U5545 ( .A(n1475), .Y(n1477) );
  INVX1 U5546 ( .A(n4757), .Y(n1459) );
endmodule


module maze_router_DW01_dec_5 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n36, n37, n38, n39, n41, n42, n43, n44, n47, n48, n49,
         n52, n53, n54, n55, n58, n59, n60, n64, n65, n70, n71, n72, n75, n76,
         n78, n79, n82, n83, n84, n88, n89, n94, n95, n96, n100, n101, n103,
         n106, n107, n108, n111, n112, n113, n118, n122, n123, n124, n127,
         n128, n129, n133, n134, n139, n140, n141, n145, n146, n148, n151,
         n152, n153, n156, n158, n163, n167, n168, n169, n172, n173, n176,
         n177, n182, n183, n187, n188, n191, n195, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351;

  XOR2X1 U12 ( .A(n298), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U21 ( .A(n297), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U28 ( .A(n296), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U44 ( .A(n295), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U53 ( .A(n294), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U60 ( .A(n293), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U76 ( .A(n292), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U92 ( .A(n328), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U101 ( .A(n340), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U108 ( .A(n335), .B(A[17]), .Y(SUM[17]) );
  XNOR2X1 U117 ( .A(n351), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U122 ( .A(n291), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U137 ( .A(n290), .B(A[13]), .Y(SUM[13]) );
  XOR2X1 U153 ( .A(n289), .B(A[11]), .Y(SUM[11]) );
  XOR2X1 U162 ( .A(n333), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U169 ( .A(n336), .B(A[9]), .Y(SUM[9]) );
  XNOR2X1 U178 ( .A(n167), .B(A[8]), .Y(SUM[8]) );
  XNOR2X1 U183 ( .A(n317), .B(A[7]), .Y(SUM[7]) );
  XNOR2X1 U191 ( .A(n288), .B(A[6]), .Y(SUM[6]) );
  XNOR2X1 U197 ( .A(n331), .B(A[5]), .Y(SUM[5]) );
  XOR2X1 U205 ( .A(n187), .B(A[4]), .Y(SUM[4]) );
  XOR2X1 U211 ( .A(n327), .B(A[3]), .Y(SUM[3]) );
  XNOR2X1 U218 ( .A(n195), .B(A[2]), .Y(SUM[2]) );
  XNOR2X1 U223 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  OR2X1 U233 ( .A(n351), .B(n310), .Y(n70) );
  AND2X1 U234 ( .A(n282), .B(n108), .Y(n107) );
  AND2X2 U235 ( .A(n278), .B(n286), .Y(n2) );
  INVX1 U236 ( .A(n2), .Y(n267) );
  OR2X2 U237 ( .A(n341), .B(n332), .Y(n37) );
  INVX1 U238 ( .A(n37), .Y(n268) );
  OR2X2 U239 ( .A(A[6]), .B(A[7]), .Y(n169) );
  INVX1 U240 ( .A(n169), .Y(n269) );
  OR2X2 U241 ( .A(A[11]), .B(A[10]), .Y(n148) );
  INVX1 U242 ( .A(n148), .Y(n270) );
  AND2X2 U243 ( .A(n270), .B(n321), .Y(n145) );
  AND2X2 U244 ( .A(n281), .B(n302), .Y(n100) );
  INVX1 U245 ( .A(n100), .Y(n271) );
  AND2X2 U246 ( .A(n303), .B(n325), .Y(n41) );
  INVX1 U247 ( .A(n41), .Y(n272) );
  AND2X2 U248 ( .A(n268), .B(n325), .Y(n36) );
  INVX1 U249 ( .A(n36), .Y(n273) );
  OR2X2 U250 ( .A(A[2]), .B(A[3]), .Y(n188) );
  INVX1 U251 ( .A(n188), .Y(n274) );
  OR2X2 U252 ( .A(n177), .B(A[6]), .Y(n173) );
  INVX1 U253 ( .A(n173), .Y(n275) );
  OR2X2 U254 ( .A(n134), .B(A[14]), .Y(n129) );
  INVX1 U255 ( .A(n129), .Y(n276) );
  OR2X2 U256 ( .A(A[23]), .B(A[22]), .Y(n79) );
  INVX1 U257 ( .A(n79), .Y(n277) );
  OR2X2 U258 ( .A(n279), .B(n322), .Y(n122) );
  INVX1 U259 ( .A(n122), .Y(n278) );
  AND2X2 U260 ( .A(n334), .B(n330), .Y(n123) );
  INVX1 U261 ( .A(n123), .Y(n279) );
  AND2X2 U262 ( .A(n269), .B(n285), .Y(n168) );
  INVX1 U263 ( .A(n168), .Y(n280) );
  OR2X2 U264 ( .A(A[17]), .B(A[16]), .Y(n113) );
  INVX1 U265 ( .A(n113), .Y(n281) );
  INVX1 U266 ( .A(n113), .Y(n282) );
  OR2X2 U267 ( .A(A[25]), .B(A[24]), .Y(n65) );
  INVX1 U268 ( .A(n65), .Y(n283) );
  OR2X2 U269 ( .A(A[9]), .B(A[8]), .Y(n158) );
  INVX1 U270 ( .A(n158), .Y(n284) );
  OR2X2 U271 ( .A(A[5]), .B(A[4]), .Y(n177) );
  INVX1 U272 ( .A(n177), .Y(n285) );
  OR2X2 U273 ( .A(n287), .B(n280), .Y(n167) );
  INVX1 U274 ( .A(n167), .Y(n286) );
  AND2X2 U275 ( .A(n274), .B(n318), .Y(n187) );
  INVX1 U276 ( .A(n187), .Y(n287) );
  AND2X2 U277 ( .A(n320), .B(n187), .Y(n176) );
  INVX1 U278 ( .A(n176), .Y(n288) );
  OR2X2 U279 ( .A(n167), .B(n305), .Y(n151) );
  INVX1 U280 ( .A(n151), .Y(n289) );
  OR2X2 U281 ( .A(n167), .B(n306), .Y(n139) );
  INVX1 U282 ( .A(n139), .Y(n290) );
  OR2X2 U283 ( .A(n167), .B(n307), .Y(n127) );
  INVX1 U284 ( .A(n127), .Y(n291) );
  OR2X1 U285 ( .A(n351), .B(n308), .Y(n94) );
  INVX1 U286 ( .A(n94), .Y(n292) );
  OR2X2 U287 ( .A(n351), .B(n309), .Y(n82) );
  INVX1 U288 ( .A(n82), .Y(n293) );
  OR2X2 U289 ( .A(n351), .B(n76), .Y(n75) );
  INVX1 U290 ( .A(n75), .Y(n294) );
  INVX1 U291 ( .A(n70), .Y(n295) );
  OR2X1 U292 ( .A(n351), .B(n311), .Y(n58) );
  INVX1 U293 ( .A(n58), .Y(n296) );
  OR2X1 U294 ( .A(n351), .B(n312), .Y(n52) );
  INVX1 U295 ( .A(n52), .Y(n297) );
  OR2X2 U296 ( .A(n351), .B(n313), .Y(n47) );
  INVX1 U297 ( .A(n47), .Y(n298) );
  OR2X2 U298 ( .A(n65), .B(A[26]), .Y(n60) );
  INVX1 U299 ( .A(n60), .Y(n299) );
  OR2X2 U300 ( .A(n342), .B(A[28]), .Y(n49) );
  INVX1 U301 ( .A(n49), .Y(n300) );
  OR2X2 U302 ( .A(n89), .B(A[22]), .Y(n84) );
  INVX1 U303 ( .A(n84), .Y(n301) );
  OR2X2 U304 ( .A(A[19]), .B(A[18]), .Y(n103) );
  INVX1 U305 ( .A(n103), .Y(n302) );
  OR2X2 U306 ( .A(n341), .B(n43), .Y(n42) );
  INVX1 U307 ( .A(n42), .Y(n303) );
  AND2X2 U308 ( .A(n339), .B(n277), .Y(n78) );
  INVX1 U309 ( .A(n78), .Y(n304) );
  AND2X2 U310 ( .A(n153), .B(n284), .Y(n152) );
  INVX1 U311 ( .A(n152), .Y(n305) );
  AND2X2 U312 ( .A(n141), .B(n146), .Y(n140) );
  INVX1 U313 ( .A(n140), .Y(n306) );
  AND2X2 U314 ( .A(n146), .B(n276), .Y(n128) );
  INVX1 U315 ( .A(n128), .Y(n307) );
  AND2X2 U316 ( .A(n96), .B(n101), .Y(n95) );
  INVX1 U317 ( .A(n95), .Y(n308) );
  AND2X2 U318 ( .A(n101), .B(n301), .Y(n83) );
  INVX1 U319 ( .A(n83), .Y(n309) );
  AND2X2 U320 ( .A(n72), .B(n325), .Y(n71) );
  INVX1 U321 ( .A(n71), .Y(n310) );
  AND2X2 U322 ( .A(n299), .B(n326), .Y(n59) );
  INVX1 U323 ( .A(n59), .Y(n311) );
  AND2X2 U324 ( .A(n54), .B(n324), .Y(n53) );
  INVX1 U325 ( .A(n53), .Y(n312) );
  AND2X2 U326 ( .A(n300), .B(n326), .Y(n48) );
  INVX1 U327 ( .A(n48), .Y(n313) );
  AND2X2 U328 ( .A(n334), .B(n146), .Y(n133) );
  INVX1 U329 ( .A(n133), .Y(n314) );
  AND2X2 U330 ( .A(n339), .B(n101), .Y(n88) );
  INVX1 U331 ( .A(n88), .Y(n315) );
  AND2X2 U332 ( .A(n319), .B(n324), .Y(n64) );
  INVX1 U333 ( .A(n64), .Y(n316) );
  AND2X2 U334 ( .A(n187), .B(n275), .Y(n172) );
  INVX1 U335 ( .A(n172), .Y(n317) );
  OR2X2 U336 ( .A(A[0]), .B(A[1]), .Y(n195) );
  INVX1 U337 ( .A(n195), .Y(n318) );
  INVX1 U338 ( .A(n65), .Y(n319) );
  INVX1 U339 ( .A(n177), .Y(n320) );
  INVX1 U340 ( .A(n158), .Y(n321) );
  OR2X2 U341 ( .A(n351), .B(n271), .Y(n349) );
  INVX1 U342 ( .A(n145), .Y(n322) );
  INVX1 U343 ( .A(n145), .Y(n323) );
  INVX1 U344 ( .A(n3), .Y(n324) );
  INVX1 U345 ( .A(n3), .Y(n325) );
  INVX1 U346 ( .A(n3), .Y(n326) );
  OR2X2 U347 ( .A(n271), .B(n304), .Y(n3) );
  OR2X2 U348 ( .A(n195), .B(A[2]), .Y(n191) );
  INVX1 U349 ( .A(n191), .Y(n327) );
  OR2X2 U350 ( .A(n351), .B(n329), .Y(n106) );
  INVX1 U351 ( .A(n106), .Y(n328) );
  INVX1 U352 ( .A(n107), .Y(n329) );
  OR2X2 U353 ( .A(A[15]), .B(A[14]), .Y(n124) );
  INVX1 U354 ( .A(n124), .Y(n330) );
  AND2X2 U355 ( .A(n183), .B(n187), .Y(n182) );
  INVX1 U356 ( .A(n182), .Y(n331) );
  AND2X2 U357 ( .A(n39), .B(n337), .Y(n38) );
  INVX1 U358 ( .A(n38), .Y(n332) );
  OR2X2 U359 ( .A(n167), .B(n158), .Y(n156) );
  INVX1 U360 ( .A(n156), .Y(n333) );
  OR2X2 U361 ( .A(A[13]), .B(A[12]), .Y(n134) );
  INVX1 U362 ( .A(n134), .Y(n334) );
  OR2X2 U363 ( .A(n351), .B(A[16]), .Y(n118) );
  INVX1 U364 ( .A(n118), .Y(n335) );
  OR2X2 U365 ( .A(n167), .B(A[8]), .Y(n163) );
  INVX1 U366 ( .A(n163), .Y(n336) );
  OR2X2 U367 ( .A(A[29]), .B(A[28]), .Y(n44) );
  INVX1 U368 ( .A(n44), .Y(n337) );
  INVX1 U369 ( .A(n44), .Y(n338) );
  OR2X2 U370 ( .A(A[21]), .B(A[20]), .Y(n89) );
  INVX1 U371 ( .A(n89), .Y(n339) );
  OR2X1 U372 ( .A(n351), .B(n112), .Y(n111) );
  INVX1 U373 ( .A(n111), .Y(n340) );
  AND2X2 U374 ( .A(n283), .B(n343), .Y(n4) );
  INVX1 U375 ( .A(n4), .Y(n341) );
  INVX1 U376 ( .A(n4), .Y(n342) );
  OR2X2 U377 ( .A(A[27]), .B(A[26]), .Y(n55) );
  INVX1 U378 ( .A(n55), .Y(n343) );
  BUFX2 U379 ( .A(n267), .Y(n351) );
  INVX1 U380 ( .A(n323), .Y(n146) );
  INVX1 U381 ( .A(n271), .Y(n101) );
  INVX1 U382 ( .A(n338), .Y(n43) );
  INVX1 U383 ( .A(n281), .Y(n112) );
  INVX1 U384 ( .A(n326), .Y(n76) );
  INVX1 U385 ( .A(n342), .Y(n54) );
  XNOR2X1 U386 ( .A(n344), .B(A[26]), .Y(SUM[26]) );
  OR2X1 U387 ( .A(n351), .B(n316), .Y(n344) );
  INVX1 U388 ( .A(A[24]), .Y(n72) );
  XNOR2X1 U389 ( .A(n345), .B(A[30]), .Y(SUM[30]) );
  OR2X1 U390 ( .A(n351), .B(n272), .Y(n345) );
  XNOR2X1 U391 ( .A(n346), .B(A[31]), .Y(SUM[31]) );
  OR2X1 U392 ( .A(n351), .B(n273), .Y(n346) );
  XNOR2X1 U393 ( .A(n347), .B(A[22]), .Y(SUM[22]) );
  OR2X1 U394 ( .A(n351), .B(n315), .Y(n347) );
  INVX1 U395 ( .A(A[20]), .Y(n96) );
  INVX1 U396 ( .A(A[18]), .Y(n108) );
  INVX1 U397 ( .A(A[10]), .Y(n153) );
  XNOR2X1 U398 ( .A(n348), .B(A[14]), .Y(SUM[14]) );
  OR2X1 U399 ( .A(n167), .B(n314), .Y(n348) );
  INVX1 U400 ( .A(A[12]), .Y(n141) );
  XNOR2X1 U401 ( .A(n349), .B(A[20]), .Y(SUM[20]) );
  XNOR2X1 U402 ( .A(n350), .B(A[12]), .Y(SUM[12]) );
  OR2X1 U403 ( .A(n167), .B(n322), .Y(n350) );
  INVX1 U404 ( .A(A[4]), .Y(n183) );
  INVX1 U405 ( .A(A[30]), .Y(n39) );
  INVX1 U406 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module maze_router_DW01_inc_6 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n23, n24, n25, n26, n29, n30, n31, n34, n35, n36, n41, n42, n45,
         n46, n47, n49, n50, n53, n54, n55, n58, n59, n60, n65, n66, n69, n70,
         n71, n72, n74, n77, n78, n81, n82, n83, n84, n89, n93, n94, n95, n98,
         n99, n100, n103, n104, n105, n110, n111, n114, n115, n117, n119, n122,
         n123, n126, n127, n128, n129, n134, n138, n139, n140, n144, n148,
         n156, n157, n158, n159, n162, n166, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322;

  XOR2X1 U6 ( .A(n264), .B(n10), .Y(SUM[30]) );
  XOR2X1 U48 ( .A(n301), .B(n45), .Y(SUM[24]) );
  XOR2X1 U76 ( .A(n303), .B(n69), .Y(SUM[20]) );
  XOR2X1 U90 ( .A(n287), .B(n81), .Y(SUM[18]) );
  XOR2X1 U129 ( .A(n294), .B(n114), .Y(SUM[12]) );
  XOR2X1 U143 ( .A(n304), .B(n126), .Y(SUM[10]) );
  XOR2X1 U180 ( .A(n157), .B(n156), .Y(SUM[4]) );
  OR2X2 U204 ( .A(n72), .B(n69), .Y(n66) );
  INVX1 U205 ( .A(n66), .Y(n238) );
  OR2X2 U206 ( .A(n72), .B(n309), .Y(n59) );
  INVX1 U207 ( .A(n59), .Y(n239) );
  OR2X2 U208 ( .A(n316), .B(n45), .Y(n42) );
  INVX1 U209 ( .A(n42), .Y(n240) );
  OR2X2 U210 ( .A(n315), .B(n279), .Y(n35) );
  INVX1 U211 ( .A(n35), .Y(n241) );
  OR2X2 U212 ( .A(n315), .B(n272), .Y(n30) );
  INVX1 U213 ( .A(n30), .Y(n242) );
  OR2X2 U214 ( .A(n316), .B(n25), .Y(n24) );
  INVX1 U215 ( .A(n24), .Y(n243) );
  OR2X2 U216 ( .A(n315), .B(n274), .Y(n19) );
  INVX1 U217 ( .A(n19), .Y(n244) );
  OR2X2 U218 ( .A(n314), .B(n275), .Y(n12) );
  INVX1 U219 ( .A(n12), .Y(n245) );
  OR2X2 U220 ( .A(n305), .B(n10), .Y(n9) );
  INVX1 U221 ( .A(n9), .Y(n246) );
  OR2X2 U222 ( .A(n316), .B(n276), .Y(n7) );
  INVX1 U223 ( .A(n7), .Y(n247) );
  OR2X2 U224 ( .A(n313), .B(n253), .Y(n139) );
  INVX1 U225 ( .A(n139), .Y(n248) );
  OR2X2 U226 ( .A(n117), .B(n114), .Y(n111) );
  INVX1 U227 ( .A(n111), .Y(n249) );
  OR2X2 U228 ( .A(n117), .B(n308), .Y(n104) );
  INVX1 U229 ( .A(n104), .Y(n250) );
  OR2X2 U230 ( .A(n117), .B(n271), .Y(n99) );
  INVX1 U231 ( .A(n99), .Y(n251) );
  AND2X2 U232 ( .A(n268), .B(n277), .Y(n93) );
  INVX1 U233 ( .A(n93), .Y(n252) );
  AND2X2 U234 ( .A(A[7]), .B(A[6]), .Y(n140) );
  INVX1 U235 ( .A(n140), .Y(n253) );
  AND2X2 U236 ( .A(n248), .B(n255), .Y(n138) );
  INVX1 U237 ( .A(n138), .Y(n254) );
  OR2X2 U238 ( .A(n257), .B(n269), .Y(n158) );
  INVX1 U239 ( .A(n158), .Y(n255) );
  INVX1 U240 ( .A(n158), .Y(n256) );
  AND2X2 U241 ( .A(A[1]), .B(A[0]), .Y(n166) );
  INVX1 U242 ( .A(n166), .Y(n257) );
  AND2X2 U243 ( .A(A[16]), .B(n2), .Y(n89) );
  INVX1 U244 ( .A(n89), .Y(n258) );
  AND2X2 U245 ( .A(n243), .B(n2), .Y(n23) );
  INVX1 U246 ( .A(n23), .Y(n259) );
  AND2X2 U247 ( .A(n244), .B(n2), .Y(n18) );
  INVX1 U248 ( .A(n18), .Y(n260) );
  AND2X2 U249 ( .A(n247), .B(n2), .Y(n6) );
  INVX1 U250 ( .A(n6), .Y(n261) );
  OR2X2 U251 ( .A(n279), .B(n273), .Y(n4) );
  INVX1 U252 ( .A(n4), .Y(n262) );
  INVX1 U253 ( .A(n4), .Y(n263) );
  AND2X2 U254 ( .A(n245), .B(n2), .Y(n11) );
  INVX1 U255 ( .A(n11), .Y(n264) );
  OR2X2 U256 ( .A(n311), .B(n270), .Y(n265) );
  OR2X2 U257 ( .A(n254), .B(n252), .Y(n319) );
  OR2X2 U258 ( .A(n312), .B(n126), .Y(n123) );
  INVX1 U259 ( .A(n123), .Y(n266) );
  OR2X2 U260 ( .A(n307), .B(n81), .Y(n78) );
  INVX1 U261 ( .A(n78), .Y(n267) );
  OR2X2 U262 ( .A(n308), .B(n290), .Y(n94) );
  INVX1 U263 ( .A(n94), .Y(n268) );
  AND2X2 U264 ( .A(A[3]), .B(A[2]), .Y(n159) );
  INVX1 U265 ( .A(n159), .Y(n269) );
  AND2X2 U266 ( .A(A[11]), .B(A[10]), .Y(n119) );
  INVX1 U267 ( .A(n119), .Y(n270) );
  AND2X2 U268 ( .A(A[14]), .B(n105), .Y(n100) );
  INVX1 U269 ( .A(n100), .Y(n271) );
  AND2X2 U270 ( .A(A[26]), .B(n36), .Y(n31) );
  INVX1 U271 ( .A(n31), .Y(n272) );
  AND2X2 U272 ( .A(A[27]), .B(A[26]), .Y(n26) );
  INVX1 U273 ( .A(n26), .Y(n273) );
  AND2X2 U274 ( .A(A[28]), .B(n262), .Y(n20) );
  INVX1 U275 ( .A(n20), .Y(n274) );
  AND2X2 U276 ( .A(n14), .B(n262), .Y(n13) );
  INVX1 U277 ( .A(n13), .Y(n275) );
  AND2X2 U278 ( .A(n246), .B(n263), .Y(n8) );
  INVX1 U279 ( .A(n8), .Y(n276) );
  INVX1 U280 ( .A(n265), .Y(n277) );
  INVX1 U281 ( .A(n265), .Y(n278) );
  INVX1 U282 ( .A(n36), .Y(n279) );
  AND2X2 U283 ( .A(A[25]), .B(A[24]), .Y(n36) );
  AND2X2 U284 ( .A(n242), .B(n2), .Y(n29) );
  INVX1 U285 ( .A(n29), .Y(n280) );
  AND2X2 U286 ( .A(n241), .B(n2), .Y(n34) );
  INVX1 U287 ( .A(n34), .Y(n281) );
  AND2X2 U288 ( .A(n240), .B(n2), .Y(n41) );
  INVX1 U289 ( .A(n41), .Y(n282) );
  AND2X2 U290 ( .A(n251), .B(n138), .Y(n98) );
  INVX1 U291 ( .A(n98), .Y(n283) );
  AND2X2 U292 ( .A(n288), .B(n2), .Y(n53) );
  INVX1 U293 ( .A(n53), .Y(n284) );
  AND2X2 U294 ( .A(n266), .B(n138), .Y(n122) );
  INVX1 U295 ( .A(n122), .Y(n285) );
  AND2X2 U296 ( .A(n267), .B(n2), .Y(n77) );
  INVX1 U297 ( .A(n77), .Y(n286) );
  AND2X2 U298 ( .A(n83), .B(n2), .Y(n82) );
  INVX1 U299 ( .A(n82), .Y(n287) );
  OR2X2 U300 ( .A(n72), .B(n289), .Y(n54) );
  INVX1 U301 ( .A(n54), .Y(n288) );
  AND2X2 U302 ( .A(A[22]), .B(n60), .Y(n55) );
  INVX1 U303 ( .A(n55), .Y(n289) );
  AND2X2 U304 ( .A(A[15]), .B(A[14]), .Y(n95) );
  INVX1 U305 ( .A(n95), .Y(n290) );
  AND2X2 U306 ( .A(A[2]), .B(n166), .Y(n162) );
  INVX1 U307 ( .A(n162), .Y(n291) );
  AND2X2 U308 ( .A(n249), .B(n138), .Y(n110) );
  INVX1 U309 ( .A(n110), .Y(n292) );
  AND2X2 U310 ( .A(n239), .B(n2), .Y(n58) );
  INVX1 U311 ( .A(n58), .Y(n293) );
  AND2X2 U312 ( .A(n277), .B(n138), .Y(n115) );
  INVX1 U313 ( .A(n115), .Y(n294) );
  OR2X2 U314 ( .A(n306), .B(n298), .Y(n71) );
  INVX1 U315 ( .A(n71), .Y(n295) );
  INVX1 U316 ( .A(n71), .Y(n296) );
  INVX1 U317 ( .A(n71), .Y(n297) );
  AND2X2 U318 ( .A(A[19]), .B(A[18]), .Y(n74) );
  INVX1 U319 ( .A(n74), .Y(n298) );
  AND2X2 U320 ( .A(A[6]), .B(n148), .Y(n144) );
  INVX1 U321 ( .A(n144), .Y(n299) );
  OR2X2 U322 ( .A(n157), .B(n299), .Y(n322) );
  AND2X2 U323 ( .A(A[8]), .B(n138), .Y(n134) );
  INVX1 U324 ( .A(n134), .Y(n300) );
  AND2X2 U325 ( .A(n47), .B(n2), .Y(n46) );
  INVX1 U326 ( .A(n46), .Y(n301) );
  AND2X2 U327 ( .A(n250), .B(n138), .Y(n103) );
  INVX1 U328 ( .A(n103), .Y(n302) );
  AND2X2 U329 ( .A(n295), .B(n2), .Y(n70) );
  INVX1 U330 ( .A(n70), .Y(n303) );
  AND2X2 U331 ( .A(n128), .B(n138), .Y(n127) );
  INVX1 U332 ( .A(n127), .Y(n304) );
  AND2X2 U333 ( .A(A[29]), .B(A[28]), .Y(n15) );
  INVX1 U334 ( .A(n15), .Y(n305) );
  AND2X2 U335 ( .A(A[17]), .B(A[16]), .Y(n84) );
  INVX1 U336 ( .A(n84), .Y(n306) );
  INVX1 U337 ( .A(n84), .Y(n307) );
  AND2X2 U338 ( .A(A[13]), .B(A[12]), .Y(n105) );
  INVX1 U339 ( .A(n105), .Y(n308) );
  AND2X2 U340 ( .A(A[21]), .B(A[20]), .Y(n60) );
  INVX1 U341 ( .A(n60), .Y(n309) );
  AND2X2 U342 ( .A(n238), .B(n2), .Y(n65) );
  INVX1 U343 ( .A(n65), .Y(n310) );
  INVX4 U344 ( .A(n319), .Y(n2) );
  AND2X2 U345 ( .A(A[9]), .B(A[8]), .Y(n129) );
  INVX1 U346 ( .A(n129), .Y(n311) );
  INVX1 U347 ( .A(n129), .Y(n312) );
  AND2X2 U348 ( .A(A[5]), .B(A[4]), .Y(n148) );
  INVX1 U349 ( .A(n148), .Y(n313) );
  OR2X2 U350 ( .A(n157), .B(n313), .Y(n321) );
  AND2X2 U351 ( .A(n317), .B(n296), .Y(n3) );
  INVX1 U352 ( .A(n3), .Y(n314) );
  INVX1 U353 ( .A(n3), .Y(n315) );
  INVX1 U354 ( .A(n3), .Y(n316) );
  OR2X2 U355 ( .A(n309), .B(n318), .Y(n49) );
  INVX1 U356 ( .A(n49), .Y(n317) );
  AND2X2 U357 ( .A(A[23]), .B(A[22]), .Y(n50) );
  INVX1 U358 ( .A(n50), .Y(n318) );
  INVX1 U359 ( .A(n305), .Y(n14) );
  INVX1 U360 ( .A(n263), .Y(n25) );
  INVX1 U361 ( .A(n256), .Y(n157) );
  INVX1 U362 ( .A(n278), .Y(n117) );
  INVX1 U363 ( .A(n297), .Y(n72) );
  INVX1 U364 ( .A(n314), .Y(n47) );
  INVX1 U365 ( .A(n312), .Y(n128) );
  INVX1 U366 ( .A(n307), .Y(n83) );
  INVX1 U367 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U368 ( .A(A[0]), .B(A[1]), .Y(SUM[1]) );
  XOR2X1 U369 ( .A(n166), .B(A[2]), .Y(SUM[2]) );
  XNOR2X1 U370 ( .A(n291), .B(A[3]), .Y(SUM[3]) );
  XNOR2X1 U371 ( .A(n320), .B(A[5]), .Y(SUM[5]) );
  OR2X1 U372 ( .A(n157), .B(n156), .Y(n320) );
  XNOR2X1 U373 ( .A(n258), .B(A[17]), .Y(SUM[17]) );
  INVX1 U374 ( .A(A[24]), .Y(n45) );
  INVX1 U375 ( .A(A[20]), .Y(n69) );
  INVX1 U376 ( .A(A[10]), .Y(n126) );
  INVX1 U377 ( .A(A[18]), .Y(n81) );
  INVX1 U378 ( .A(A[12]), .Y(n114) );
  INVX1 U379 ( .A(A[30]), .Y(n10) );
  XNOR2X1 U380 ( .A(n292), .B(A[13]), .Y(SUM[13]) );
  XNOR2X1 U381 ( .A(n286), .B(A[19]), .Y(SUM[19]) );
  XNOR2X1 U382 ( .A(n310), .B(A[21]), .Y(SUM[21]) );
  XNOR2X1 U383 ( .A(n293), .B(A[22]), .Y(SUM[22]) );
  XNOR2X1 U384 ( .A(n284), .B(A[23]), .Y(SUM[23]) );
  XNOR2X1 U385 ( .A(n282), .B(A[25]), .Y(SUM[25]) );
  XNOR2X1 U386 ( .A(n281), .B(A[26]), .Y(SUM[26]) );
  XNOR2X1 U387 ( .A(n280), .B(A[27]), .Y(SUM[27]) );
  XNOR2X1 U388 ( .A(n259), .B(A[28]), .Y(SUM[28]) );
  XNOR2X1 U389 ( .A(n260), .B(A[29]), .Y(SUM[29]) );
  XNOR2X1 U390 ( .A(n261), .B(A[31]), .Y(SUM[31]) );
  XNOR2X1 U391 ( .A(n321), .B(A[6]), .Y(SUM[6]) );
  XNOR2X1 U392 ( .A(n322), .B(A[7]), .Y(SUM[7]) );
  XOR2X1 U393 ( .A(n138), .B(A[8]), .Y(SUM[8]) );
  XNOR2X1 U394 ( .A(n300), .B(A[9]), .Y(SUM[9]) );
  XNOR2X1 U395 ( .A(n285), .B(A[11]), .Y(SUM[11]) );
  XNOR2X1 U396 ( .A(n302), .B(A[14]), .Y(SUM[14]) );
  XNOR2X1 U397 ( .A(n283), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U398 ( .A(n2), .B(A[16]), .Y(SUM[16]) );
  INVX1 U399 ( .A(A[4]), .Y(n156) );
endmodule


module maze_router_DW01_inc_7 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n23, n24, n25, n26, n29, n30, n31, n34, n35, n36, n41, n42, n45,
         n46, n47, n49, n50, n53, n54, n55, n58, n59, n60, n65, n66, n69, n70,
         n71, n72, n74, n77, n78, n81, n82, n84, n89, n93, n94, n95, n98, n99,
         n100, n103, n104, n105, n110, n111, n114, n115, n116, n119, n122,
         n123, n126, n127, n129, n134, n138, n139, n140, n142, n143, n144,
         n148, n156, n157, n158, n159, n162, n166, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;

  XOR2X1 U6 ( .A(n284), .B(n10), .Y(SUM[30]) );
  XOR2X1 U48 ( .A(n283), .B(n45), .Y(SUM[24]) );
  XOR2X1 U76 ( .A(n282), .B(n69), .Y(SUM[20]) );
  XOR2X1 U90 ( .A(n281), .B(n81), .Y(SUM[18]) );
  XOR2X1 U129 ( .A(n280), .B(n114), .Y(SUM[12]) );
  XOR2X1 U143 ( .A(n279), .B(n126), .Y(SUM[10]) );
  XNOR2X1 U161 ( .A(n306), .B(n142), .Y(SUM[7]) );
  XOR2X1 U180 ( .A(n157), .B(n156), .Y(SUM[4]) );
  OR2X2 U204 ( .A(n116), .B(n114), .Y(n111) );
  INVX1 U205 ( .A(n111), .Y(n238) );
  OR2X2 U206 ( .A(n116), .B(n312), .Y(n104) );
  INVX1 U207 ( .A(n104), .Y(n239) );
  OR2X2 U208 ( .A(n116), .B(n308), .Y(n99) );
  INVX1 U209 ( .A(n99), .Y(n240) );
  OR2X2 U210 ( .A(n72), .B(n69), .Y(n66) );
  INVX1 U211 ( .A(n66), .Y(n241) );
  OR2X2 U212 ( .A(n72), .B(n315), .Y(n59) );
  INVX1 U213 ( .A(n59), .Y(n242) );
  OR2X2 U214 ( .A(n72), .B(n311), .Y(n54) );
  INVX1 U215 ( .A(n54), .Y(n243) );
  OR2X2 U216 ( .A(n304), .B(n45), .Y(n42) );
  INVX1 U217 ( .A(n42), .Y(n244) );
  OR2X2 U218 ( .A(n304), .B(n253), .Y(n35) );
  INVX1 U219 ( .A(n35), .Y(n245) );
  OR2X2 U220 ( .A(n303), .B(n291), .Y(n30) );
  INVX1 U221 ( .A(n30), .Y(n246) );
  OR2X2 U222 ( .A(n304), .B(n292), .Y(n19) );
  INVX1 U223 ( .A(n19), .Y(n247) );
  OR2X2 U224 ( .A(n304), .B(n293), .Y(n12) );
  INVX1 U225 ( .A(n12), .Y(n248) );
  OR2X2 U226 ( .A(n304), .B(n294), .Y(n7) );
  INVX1 U227 ( .A(n7), .Y(n249) );
  AND2X2 U228 ( .A(A[11]), .B(A[10]), .Y(n119) );
  INVX1 U229 ( .A(n119), .Y(n250) );
  OR2X2 U230 ( .A(n262), .B(n250), .Y(n116) );
  AND2X2 U231 ( .A(n256), .B(n296), .Y(n93) );
  INVX1 U232 ( .A(n93), .Y(n251) );
  OR2X2 U233 ( .A(n263), .B(n290), .Y(n71) );
  OR2X2 U234 ( .A(n315), .B(n258), .Y(n49) );
  INVX1 U235 ( .A(n49), .Y(n252) );
  AND2X2 U236 ( .A(n252), .B(n297), .Y(n3) );
  AND2X2 U237 ( .A(A[25]), .B(A[24]), .Y(n36) );
  INVX1 U238 ( .A(n36), .Y(n253) );
  OR2X2 U239 ( .A(n253), .B(n259), .Y(n4) );
  OR2X2 U240 ( .A(n314), .B(n10), .Y(n9) );
  INVX1 U241 ( .A(n9), .Y(n254) );
  OR2X2 U242 ( .A(n313), .B(n288), .Y(n139) );
  INVX1 U243 ( .A(n139), .Y(n255) );
  OR2X2 U244 ( .A(n312), .B(n289), .Y(n94) );
  INVX1 U245 ( .A(n94), .Y(n256) );
  AND2X2 U246 ( .A(A[3]), .B(A[2]), .Y(n159) );
  INVX1 U247 ( .A(n159), .Y(n257) );
  AND2X2 U248 ( .A(A[23]), .B(A[22]), .Y(n50) );
  INVX1 U249 ( .A(n50), .Y(n258) );
  AND2X2 U250 ( .A(A[27]), .B(A[26]), .Y(n26) );
  INVX1 U251 ( .A(n26), .Y(n259) );
  OR2X2 U252 ( .A(n257), .B(n295), .Y(n158) );
  INVX1 U253 ( .A(n158), .Y(n260) );
  INVX1 U254 ( .A(n158), .Y(n261) );
  AND2X2 U255 ( .A(A[9]), .B(A[8]), .Y(n129) );
  INVX1 U256 ( .A(n129), .Y(n262) );
  AND2X2 U257 ( .A(A[17]), .B(A[16]), .Y(n84) );
  INVX1 U258 ( .A(n84), .Y(n263) );
  AND2X2 U259 ( .A(n260), .B(n255), .Y(n138) );
  INVX1 U260 ( .A(n138), .Y(n264) );
  AND2X2 U261 ( .A(n286), .B(n138), .Y(n122) );
  INVX1 U262 ( .A(n122), .Y(n265) );
  AND2X2 U263 ( .A(n138), .B(n238), .Y(n110) );
  INVX1 U264 ( .A(n110), .Y(n266) );
  AND2X2 U265 ( .A(n138), .B(n239), .Y(n103) );
  INVX1 U266 ( .A(n103), .Y(n267) );
  AND2X2 U267 ( .A(n138), .B(n240), .Y(n98) );
  INVX1 U268 ( .A(n98), .Y(n268) );
  AND2X2 U269 ( .A(n287), .B(n2), .Y(n77) );
  INVX1 U270 ( .A(n77), .Y(n269) );
  AND2X2 U271 ( .A(n241), .B(n2), .Y(n65) );
  INVX1 U272 ( .A(n65), .Y(n270) );
  AND2X2 U273 ( .A(n242), .B(n2), .Y(n58) );
  INVX1 U274 ( .A(n58), .Y(n271) );
  AND2X2 U275 ( .A(n243), .B(n2), .Y(n53) );
  INVX1 U276 ( .A(n53), .Y(n272) );
  AND2X2 U277 ( .A(n2), .B(n244), .Y(n41) );
  INVX1 U278 ( .A(n41), .Y(n273) );
  AND2X2 U279 ( .A(n2), .B(n245), .Y(n34) );
  INVX1 U280 ( .A(n34), .Y(n274) );
  AND2X2 U281 ( .A(n2), .B(n246), .Y(n29) );
  INVX1 U282 ( .A(n29), .Y(n275) );
  AND2X2 U283 ( .A(n2), .B(n285), .Y(n23) );
  INVX1 U284 ( .A(n23), .Y(n276) );
  AND2X2 U285 ( .A(n2), .B(n247), .Y(n18) );
  INVX1 U286 ( .A(n18), .Y(n277) );
  AND2X2 U287 ( .A(n2), .B(n249), .Y(n6) );
  INVX1 U288 ( .A(n6), .Y(n278) );
  AND2X2 U289 ( .A(n129), .B(n138), .Y(n127) );
  INVX1 U290 ( .A(n127), .Y(n279) );
  AND2X2 U291 ( .A(n296), .B(n138), .Y(n115) );
  INVX1 U292 ( .A(n115), .Y(n280) );
  AND2X2 U293 ( .A(n84), .B(n2), .Y(n82) );
  INVX1 U294 ( .A(n82), .Y(n281) );
  AND2X2 U295 ( .A(n297), .B(n2), .Y(n70) );
  INVX1 U296 ( .A(n70), .Y(n282) );
  AND2X2 U297 ( .A(n47), .B(n2), .Y(n46) );
  INVX1 U298 ( .A(n46), .Y(n283) );
  AND2X2 U299 ( .A(n2), .B(n248), .Y(n11) );
  INVX1 U300 ( .A(n11), .Y(n284) );
  OR2X2 U301 ( .A(n303), .B(n25), .Y(n24) );
  INVX1 U302 ( .A(n24), .Y(n285) );
  OR2X2 U303 ( .A(n299), .B(n126), .Y(n123) );
  INVX1 U304 ( .A(n123), .Y(n286) );
  OR2X2 U305 ( .A(n300), .B(n81), .Y(n78) );
  INVX1 U306 ( .A(n78), .Y(n287) );
  AND2X2 U307 ( .A(A[7]), .B(A[6]), .Y(n140) );
  INVX1 U308 ( .A(n140), .Y(n288) );
  AND2X2 U309 ( .A(A[15]), .B(A[14]), .Y(n95) );
  INVX1 U310 ( .A(n95), .Y(n289) );
  AND2X2 U311 ( .A(A[19]), .B(A[18]), .Y(n74) );
  INVX1 U312 ( .A(n74), .Y(n290) );
  AND2X2 U313 ( .A(A[26]), .B(n36), .Y(n31) );
  INVX1 U314 ( .A(n31), .Y(n291) );
  AND2X2 U315 ( .A(A[28]), .B(n301), .Y(n20) );
  INVX1 U316 ( .A(n20), .Y(n292) );
  AND2X2 U317 ( .A(n14), .B(n302), .Y(n13) );
  INVX1 U318 ( .A(n13), .Y(n293) );
  AND2X2 U319 ( .A(n254), .B(n302), .Y(n8) );
  INVX1 U320 ( .A(n8), .Y(n294) );
  AND2X2 U321 ( .A(A[0]), .B(A[1]), .Y(n166) );
  INVX1 U322 ( .A(n166), .Y(n295) );
  INVX1 U323 ( .A(n116), .Y(n296) );
  INVX1 U324 ( .A(n71), .Y(n297) );
  INVX1 U325 ( .A(n71), .Y(n298) );
  INVX1 U326 ( .A(n129), .Y(n299) );
  INVX1 U327 ( .A(n84), .Y(n300) );
  INVX1 U328 ( .A(n4), .Y(n301) );
  INVX1 U329 ( .A(n4), .Y(n302) );
  INVX1 U330 ( .A(n3), .Y(n303) );
  INVX1 U331 ( .A(n3), .Y(n304) );
  AND2X2 U332 ( .A(A[2]), .B(n166), .Y(n162) );
  INVX1 U333 ( .A(n162), .Y(n305) );
  OR2X2 U334 ( .A(n157), .B(n307), .Y(n143) );
  INVX1 U335 ( .A(n143), .Y(n306) );
  AND2X2 U336 ( .A(A[6]), .B(n148), .Y(n144) );
  INVX1 U337 ( .A(n144), .Y(n307) );
  AND2X2 U338 ( .A(A[14]), .B(n105), .Y(n100) );
  INVX1 U339 ( .A(n100), .Y(n308) );
  AND2X2 U340 ( .A(A[16]), .B(n2), .Y(n89) );
  INVX1 U341 ( .A(n89), .Y(n309) );
  INVX4 U342 ( .A(n316), .Y(n2) );
  AND2X2 U343 ( .A(A[8]), .B(n138), .Y(n134) );
  INVX1 U344 ( .A(n134), .Y(n310) );
  AND2X2 U345 ( .A(A[22]), .B(n60), .Y(n55) );
  INVX1 U346 ( .A(n55), .Y(n311) );
  AND2X2 U347 ( .A(A[13]), .B(A[12]), .Y(n105) );
  INVX1 U348 ( .A(n105), .Y(n312) );
  AND2X2 U349 ( .A(A[4]), .B(A[5]), .Y(n148) );
  INVX1 U350 ( .A(n148), .Y(n313) );
  OR2X2 U351 ( .A(n157), .B(n313), .Y(n318) );
  AND2X2 U352 ( .A(A[29]), .B(A[28]), .Y(n15) );
  INVX1 U353 ( .A(n15), .Y(n314) );
  AND2X2 U354 ( .A(A[21]), .B(A[20]), .Y(n60) );
  INVX1 U355 ( .A(n60), .Y(n315) );
  OR2X1 U356 ( .A(n251), .B(n264), .Y(n316) );
  INVX1 U357 ( .A(n303), .Y(n47) );
  INVX1 U358 ( .A(n261), .Y(n157) );
  INVX1 U359 ( .A(n298), .Y(n72) );
  INVX1 U360 ( .A(n301), .Y(n25) );
  INVX1 U361 ( .A(n314), .Y(n14) );
  XNOR2X1 U362 ( .A(n268), .B(A[15]), .Y(SUM[15]) );
  XNOR2X1 U363 ( .A(n274), .B(A[26]), .Y(SUM[26]) );
  XNOR2X1 U364 ( .A(n278), .B(A[31]), .Y(SUM[31]) );
  XNOR2X1 U365 ( .A(n275), .B(A[27]), .Y(SUM[27]) );
  XNOR2X1 U366 ( .A(n273), .B(A[25]), .Y(SUM[25]) );
  XNOR2X1 U367 ( .A(n272), .B(A[23]), .Y(SUM[23]) );
  XNOR2X1 U368 ( .A(n270), .B(A[21]), .Y(SUM[21]) );
  XNOR2X1 U369 ( .A(n309), .B(A[17]), .Y(SUM[17]) );
  XNOR2X1 U370 ( .A(n269), .B(A[19]), .Y(SUM[19]) );
  XNOR2X1 U371 ( .A(n277), .B(A[29]), .Y(SUM[29]) );
  XNOR2X1 U372 ( .A(n265), .B(A[11]), .Y(SUM[11]) );
  XNOR2X1 U373 ( .A(n310), .B(A[9]), .Y(SUM[9]) );
  XNOR2X1 U374 ( .A(n266), .B(A[13]), .Y(SUM[13]) );
  XNOR2X1 U375 ( .A(n305), .B(A[3]), .Y(SUM[3]) );
  XNOR2X1 U376 ( .A(n276), .B(A[28]), .Y(SUM[28]) );
  XNOR2X1 U377 ( .A(n271), .B(A[22]), .Y(SUM[22]) );
  XNOR2X1 U378 ( .A(n267), .B(A[14]), .Y(SUM[14]) );
  INVX1 U379 ( .A(A[7]), .Y(n142) );
  XNOR2X1 U380 ( .A(n317), .B(A[5]), .Y(SUM[5]) );
  OR2X1 U381 ( .A(n157), .B(n156), .Y(n317) );
  XOR2X1 U382 ( .A(n138), .B(A[8]), .Y(SUM[8]) );
  XOR2X1 U383 ( .A(n2), .B(A[16]), .Y(SUM[16]) );
  XNOR2X1 U384 ( .A(n318), .B(A[6]), .Y(SUM[6]) );
  XOR2X1 U385 ( .A(n166), .B(A[2]), .Y(SUM[2]) );
  XOR2X1 U386 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  INVX1 U387 ( .A(A[0]), .Y(SUM[0]) );
  INVX1 U388 ( .A(A[4]), .Y(n156) );
  INVX1 U389 ( .A(A[24]), .Y(n45) );
  INVX1 U390 ( .A(A[18]), .Y(n81) );
  INVX1 U391 ( .A(A[20]), .Y(n69) );
  INVX1 U392 ( .A(A[12]), .Y(n114) );
  INVX1 U393 ( .A(A[10]), .Y(n126) );
  INVX1 U394 ( .A(A[30]), .Y(n10) );
endmodule


module maze_router_DW_leftsh_3 ( A, SH, B );
  input [179:0] A;
  input [31:0] SH;
  output [179:0] B;
  wire   n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n874, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1784, n1791, n1792,
         n1793, n1794, n1801, n1802, n1803, n1804, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;

  AND2X1 U50 ( .A(n355), .B(n2384), .Y(B[161]) );
  MUX2X1 U374 ( .B(n681), .A(n617), .S(n2406), .Y(n373) );
  MUX2X1 U375 ( .B(n680), .A(n616), .S(n2406), .Y(n372) );
  MUX2X1 U376 ( .B(n679), .A(n615), .S(n2406), .Y(n371) );
  MUX2X1 U377 ( .B(n678), .A(n614), .S(n2406), .Y(n370) );
  MUX2X1 U378 ( .B(n677), .A(n613), .S(n2406), .Y(n369) );
  MUX2X1 U379 ( .B(n676), .A(n612), .S(n2406), .Y(n368) );
  MUX2X1 U380 ( .B(n675), .A(n611), .S(n2406), .Y(n367) );
  MUX2X1 U381 ( .B(n674), .A(n610), .S(n2406), .Y(n366) );
  MUX2X1 U382 ( .B(n673), .A(n609), .S(n2406), .Y(n365) );
  MUX2X1 U383 ( .B(n672), .A(n608), .S(n2406), .Y(n364) );
  MUX2X1 U384 ( .B(n671), .A(n607), .S(n2406), .Y(n363) );
  MUX2X1 U385 ( .B(n670), .A(n606), .S(n2406), .Y(n362) );
  MUX2X1 U386 ( .B(n669), .A(n605), .S(n2407), .Y(n361) );
  MUX2X1 U387 ( .B(n668), .A(n604), .S(n2407), .Y(n360) );
  MUX2X1 U388 ( .B(n667), .A(n603), .S(n2407), .Y(n359) );
  MUX2X1 U389 ( .B(n666), .A(n602), .S(n2407), .Y(n358) );
  MUX2X1 U390 ( .B(n665), .A(n601), .S(n2407), .Y(n357) );
  MUX2X1 U391 ( .B(n664), .A(n600), .S(n2407), .Y(n356) );
  MUX2X1 U392 ( .B(n663), .A(n599), .S(n2407), .Y(n355) );
  MUX2X1 U393 ( .B(n662), .A(n598), .S(n2407), .Y(n354) );
  MUX2X1 U394 ( .B(n661), .A(n597), .S(n2407), .Y(n353) );
  MUX2X1 U395 ( .B(n660), .A(n596), .S(n2407), .Y(n352) );
  MUX2X1 U396 ( .B(n659), .A(n595), .S(n2407), .Y(n351) );
  MUX2X1 U397 ( .B(n658), .A(n594), .S(n2407), .Y(n350) );
  MUX2X1 U398 ( .B(n657), .A(n593), .S(n2408), .Y(n349) );
  MUX2X1 U399 ( .B(n656), .A(n592), .S(n2408), .Y(n348) );
  MUX2X1 U400 ( .B(n655), .A(n591), .S(n2408), .Y(n347) );
  MUX2X1 U401 ( .B(n654), .A(n590), .S(n2408), .Y(n346) );
  MUX2X1 U402 ( .B(n653), .A(n589), .S(n2408), .Y(n345) );
  MUX2X1 U403 ( .B(n652), .A(n588), .S(n2408), .Y(n344) );
  MUX2X1 U404 ( .B(n651), .A(n587), .S(n2408), .Y(n343) );
  MUX2X1 U405 ( .B(n650), .A(n586), .S(n2408), .Y(n342) );
  MUX2X1 U406 ( .B(n649), .A(n585), .S(n2408), .Y(n341) );
  MUX2X1 U407 ( .B(n648), .A(n584), .S(n2408), .Y(n340) );
  MUX2X1 U408 ( .B(n647), .A(n583), .S(n2408), .Y(n339) );
  MUX2X1 U409 ( .B(n646), .A(n582), .S(n2408), .Y(n338) );
  MUX2X1 U410 ( .B(n645), .A(n581), .S(n2409), .Y(n337) );
  MUX2X1 U411 ( .B(n644), .A(n580), .S(n2409), .Y(n336) );
  MUX2X1 U412 ( .B(n643), .A(n579), .S(n2409), .Y(n335) );
  MUX2X1 U413 ( .B(n642), .A(n578), .S(n2409), .Y(n334) );
  MUX2X1 U414 ( .B(n641), .A(n577), .S(n2409), .Y(n333) );
  MUX2X1 U415 ( .B(n640), .A(n576), .S(n2409), .Y(n332) );
  MUX2X1 U416 ( .B(n639), .A(n575), .S(n2409), .Y(n331) );
  MUX2X1 U417 ( .B(n638), .A(n574), .S(n2409), .Y(n330) );
  MUX2X1 U418 ( .B(n637), .A(n573), .S(n2409), .Y(n329) );
  MUX2X1 U419 ( .B(n636), .A(n572), .S(n2409), .Y(n328) );
  MUX2X1 U420 ( .B(n635), .A(n571), .S(n2409), .Y(n327) );
  MUX2X1 U421 ( .B(n634), .A(n570), .S(n2409), .Y(n326) );
  MUX2X1 U422 ( .B(n633), .A(n569), .S(n2410), .Y(n325) );
  MUX2X1 U423 ( .B(n632), .A(n568), .S(n2410), .Y(n324) );
  MUX2X1 U424 ( .B(n631), .A(n567), .S(n2410), .Y(n323) );
  MUX2X1 U425 ( .B(n630), .A(n566), .S(n2410), .Y(n322) );
  MUX2X1 U426 ( .B(n629), .A(n565), .S(n2410), .Y(n321) );
  MUX2X1 U427 ( .B(n628), .A(n564), .S(n2410), .Y(n320) );
  MUX2X1 U428 ( .B(n627), .A(n563), .S(n2410), .Y(n319) );
  MUX2X1 U429 ( .B(n626), .A(n562), .S(n2410), .Y(n318) );
  MUX2X1 U430 ( .B(n625), .A(n561), .S(n2410), .Y(n317) );
  MUX2X1 U431 ( .B(n624), .A(n560), .S(n2410), .Y(n316) );
  MUX2X1 U432 ( .B(n623), .A(n559), .S(n2410), .Y(n315) );
  MUX2X1 U433 ( .B(n622), .A(n558), .S(n2410), .Y(n314) );
  MUX2X1 U434 ( .B(n621), .A(n557), .S(n2411), .Y(n313) );
  MUX2X1 U435 ( .B(n620), .A(n556), .S(n2411), .Y(n312) );
  MUX2X1 U436 ( .B(n619), .A(n555), .S(n2411), .Y(n311) );
  MUX2X1 U437 ( .B(n618), .A(n554), .S(n2411), .Y(n310) );
  MUX2X1 U438 ( .B(n617), .A(n553), .S(n2411), .Y(n309) );
  MUX2X1 U439 ( .B(n616), .A(n552), .S(n2411), .Y(n308) );
  MUX2X1 U440 ( .B(n615), .A(n551), .S(n2411), .Y(n307) );
  MUX2X1 U441 ( .B(n614), .A(n550), .S(n2411), .Y(n306) );
  MUX2X1 U442 ( .B(n613), .A(n549), .S(n2411), .Y(n305) );
  MUX2X1 U443 ( .B(n612), .A(n548), .S(n2411), .Y(n304) );
  MUX2X1 U444 ( .B(n611), .A(n547), .S(n2411), .Y(n303) );
  MUX2X1 U445 ( .B(n610), .A(n546), .S(n2411), .Y(n302) );
  MUX2X1 U446 ( .B(n609), .A(n545), .S(n2412), .Y(n301) );
  MUX2X1 U447 ( .B(n608), .A(n544), .S(n2412), .Y(n300) );
  MUX2X1 U448 ( .B(n607), .A(n543), .S(n2412), .Y(n299) );
  MUX2X1 U449 ( .B(n606), .A(n542), .S(n2412), .Y(n298) );
  MUX2X1 U450 ( .B(n605), .A(n541), .S(n2412), .Y(n297) );
  MUX2X1 U451 ( .B(n604), .A(n540), .S(n2412), .Y(n296) );
  MUX2X1 U452 ( .B(n603), .A(n539), .S(n2412), .Y(n295) );
  MUX2X1 U453 ( .B(n602), .A(n538), .S(n2412), .Y(n294) );
  MUX2X1 U454 ( .B(n601), .A(n537), .S(n2412), .Y(n293) );
  MUX2X1 U455 ( .B(n600), .A(n536), .S(n2412), .Y(n292) );
  MUX2X1 U456 ( .B(n599), .A(n535), .S(n2412), .Y(n291) );
  MUX2X1 U457 ( .B(n598), .A(n534), .S(n2412), .Y(n290) );
  MUX2X1 U458 ( .B(n597), .A(n533), .S(n2413), .Y(n289) );
  MUX2X1 U459 ( .B(n596), .A(n532), .S(n2413), .Y(n288) );
  MUX2X1 U460 ( .B(n595), .A(n531), .S(n2413), .Y(n287) );
  MUX2X1 U461 ( .B(n594), .A(n530), .S(n2413), .Y(n286) );
  MUX2X1 U462 ( .B(n593), .A(n529), .S(n2413), .Y(n285) );
  MUX2X1 U463 ( .B(n592), .A(n528), .S(n2413), .Y(n284) );
  MUX2X1 U464 ( .B(n591), .A(n527), .S(n2413), .Y(n283) );
  MUX2X1 U465 ( .B(n590), .A(n526), .S(n2413), .Y(n282) );
  MUX2X1 U466 ( .B(n589), .A(n525), .S(n2413), .Y(n281) );
  MUX2X1 U467 ( .B(n588), .A(n524), .S(n2413), .Y(n280) );
  MUX2X1 U468 ( .B(n587), .A(n523), .S(n2413), .Y(n279) );
  MUX2X1 U469 ( .B(n586), .A(n522), .S(n2413), .Y(n278) );
  MUX2X1 U470 ( .B(n585), .A(n521), .S(n2414), .Y(n277) );
  MUX2X1 U471 ( .B(n584), .A(n520), .S(n2414), .Y(n276) );
  MUX2X1 U472 ( .B(n583), .A(n519), .S(n2414), .Y(n275) );
  MUX2X1 U473 ( .B(n582), .A(n518), .S(n2414), .Y(n274) );
  MUX2X1 U474 ( .B(n581), .A(n517), .S(n2414), .Y(n273) );
  MUX2X1 U475 ( .B(n580), .A(n516), .S(n2414), .Y(n272) );
  MUX2X1 U476 ( .B(n579), .A(n515), .S(n2414), .Y(n271) );
  MUX2X1 U477 ( .B(n578), .A(n514), .S(n2414), .Y(n270) );
  MUX2X1 U478 ( .B(n577), .A(n513), .S(n2414), .Y(n269) );
  MUX2X1 U479 ( .B(n576), .A(n512), .S(n2414), .Y(n268) );
  MUX2X1 U480 ( .B(n575), .A(n511), .S(n2414), .Y(n267) );
  MUX2X1 U481 ( .B(n574), .A(n510), .S(n2414), .Y(n266) );
  MUX2X1 U482 ( .B(n573), .A(n509), .S(n2415), .Y(n265) );
  MUX2X1 U483 ( .B(n572), .A(n508), .S(n2415), .Y(n264) );
  MUX2X1 U484 ( .B(n571), .A(n507), .S(n2415), .Y(n263) );
  MUX2X1 U485 ( .B(n570), .A(n506), .S(n2415), .Y(n262) );
  MUX2X1 U486 ( .B(n569), .A(n505), .S(n2415), .Y(n261) );
  MUX2X1 U487 ( .B(n568), .A(n504), .S(n2415), .Y(n260) );
  MUX2X1 U488 ( .B(n567), .A(n503), .S(n2415), .Y(n259) );
  MUX2X1 U489 ( .B(n566), .A(n502), .S(n2415), .Y(n258) );
  MUX2X1 U554 ( .B(n861), .A(n733), .S(n2389), .Y(n681) );
  MUX2X1 U555 ( .B(n860), .A(n732), .S(n2389), .Y(n680) );
  MUX2X1 U556 ( .B(n859), .A(n731), .S(n2389), .Y(n679) );
  MUX2X1 U557 ( .B(n858), .A(n730), .S(n2389), .Y(n678) );
  MUX2X1 U558 ( .B(n857), .A(n729), .S(n2389), .Y(n677) );
  MUX2X1 U559 ( .B(n856), .A(n728), .S(n2389), .Y(n676) );
  MUX2X1 U560 ( .B(n855), .A(n727), .S(n2389), .Y(n675) );
  MUX2X1 U561 ( .B(n854), .A(n726), .S(n2389), .Y(n674) );
  MUX2X1 U562 ( .B(n853), .A(n725), .S(n2389), .Y(n673) );
  MUX2X1 U563 ( .B(n852), .A(n724), .S(n2389), .Y(n672) );
  MUX2X1 U564 ( .B(n851), .A(n2332), .S(n2389), .Y(n671) );
  MUX2X1 U565 ( .B(n850), .A(n722), .S(n2389), .Y(n670) );
  MUX2X1 U566 ( .B(n849), .A(n721), .S(n2390), .Y(n669) );
  MUX2X1 U567 ( .B(n848), .A(n720), .S(n2390), .Y(n668) );
  MUX2X1 U568 ( .B(n847), .A(n719), .S(n2390), .Y(n667) );
  MUX2X1 U569 ( .B(n846), .A(n718), .S(n2390), .Y(n666) );
  MUX2X1 U570 ( .B(n845), .A(n717), .S(n2390), .Y(n665) );
  MUX2X1 U571 ( .B(n844), .A(n716), .S(n2390), .Y(n664) );
  MUX2X1 U572 ( .B(n843), .A(n715), .S(n2390), .Y(n663) );
  MUX2X1 U573 ( .B(n842), .A(n714), .S(n2390), .Y(n662) );
  MUX2X1 U574 ( .B(n841), .A(n2342), .S(n2390), .Y(n661) );
  MUX2X1 U575 ( .B(n840), .A(n2355), .S(n2390), .Y(n660) );
  MUX2X1 U576 ( .B(n839), .A(n2351), .S(n2390), .Y(n659) );
  MUX2X1 U577 ( .B(n838), .A(n2360), .S(n2390), .Y(n658) );
  MUX2X1 U578 ( .B(n837), .A(n2314), .S(n2391), .Y(n657) );
  MUX2X1 U579 ( .B(n836), .A(n2340), .S(n2391), .Y(n656) );
  MUX2X1 U580 ( .B(n835), .A(n2344), .S(n2391), .Y(n655) );
  MUX2X1 U581 ( .B(n834), .A(n2365), .S(n2391), .Y(n654) );
  MUX2X1 U582 ( .B(n833), .A(n2348), .S(n2391), .Y(n653) );
  MUX2X1 U583 ( .B(n832), .A(n2369), .S(n2391), .Y(n652) );
  MUX2X1 U584 ( .B(n831), .A(n2338), .S(n2391), .Y(n651) );
  MUX2X1 U585 ( .B(n830), .A(n2357), .S(n2391), .Y(n650) );
  MUX2X1 U586 ( .B(n829), .A(n2230), .S(n2391), .Y(n649) );
  MUX2X1 U587 ( .B(n828), .A(n2353), .S(n2391), .Y(n648) );
  MUX2X1 U588 ( .B(n827), .A(n2341), .S(n2391), .Y(n647) );
  MUX2X1 U589 ( .B(n826), .A(n2349), .S(n2397), .Y(n646) );
  MUX2X1 U590 ( .B(n825), .A(n2345), .S(n2392), .Y(n645) );
  MUX2X1 U591 ( .B(n824), .A(n2354), .S(n2392), .Y(n644) );
  MUX2X1 U592 ( .B(n823), .A(n2356), .S(n2392), .Y(n643) );
  MUX2X1 U593 ( .B(n822), .A(n2362), .S(n2392), .Y(n642) );
  MUX2X1 U594 ( .B(n821), .A(n2313), .S(n2392), .Y(n641) );
  MUX2X1 U595 ( .B(n820), .A(n2312), .S(n2392), .Y(n640) );
  MUX2X1 U596 ( .B(n819), .A(n2352), .S(n2392), .Y(n639) );
  MUX2X1 U597 ( .B(n818), .A(n2370), .S(n2392), .Y(n638) );
  MUX2X1 U598 ( .B(n817), .A(n2339), .S(n2392), .Y(n637) );
  MUX2X1 U599 ( .B(n816), .A(n2359), .S(n2392), .Y(n636) );
  MUX2X1 U600 ( .B(n815), .A(n2343), .S(n2392), .Y(n635) );
  MUX2X1 U601 ( .B(n814), .A(n2366), .S(n2392), .Y(n634) );
  MUX2X1 U602 ( .B(n813), .A(n2311), .S(n2393), .Y(n633) );
  MUX2X1 U603 ( .B(n812), .A(n2310), .S(n2393), .Y(n632) );
  MUX2X1 U604 ( .B(n811), .A(n2309), .S(n2393), .Y(n631) );
  MUX2X1 U605 ( .B(n810), .A(n2227), .S(n2393), .Y(n630) );
  OR2X1 U606 ( .A(n2393), .B(n374), .Y(n629) );
  OR2X1 U608 ( .A(n2393), .B(n375), .Y(n628) );
  OR2X1 U610 ( .A(n2393), .B(n376), .Y(n627) );
  OR2X1 U612 ( .A(n2393), .B(n377), .Y(n626) );
  OR2X1 U614 ( .A(n2393), .B(n378), .Y(n625) );
  OR2X1 U616 ( .A(n2393), .B(n379), .Y(n624) );
  OR2X1 U618 ( .A(n2393), .B(n380), .Y(n623) );
  OR2X1 U620 ( .A(n2393), .B(n381), .Y(n622) );
  OR2X1 U622 ( .A(n2393), .B(n382), .Y(n621) );
  OR2X1 U624 ( .A(n2393), .B(n383), .Y(n620) );
  OR2X1 U626 ( .A(n2393), .B(n384), .Y(n619) );
  OR2X1 U628 ( .A(n2393), .B(n385), .Y(n618) );
  OR2X1 U630 ( .A(n2393), .B(n386), .Y(n617) );
  OR2X1 U632 ( .A(n2393), .B(n387), .Y(n616) );
  OR2X1 U634 ( .A(n2394), .B(n388), .Y(n615) );
  OR2X1 U636 ( .A(n2394), .B(n389), .Y(n614) );
  OR2X1 U638 ( .A(n2394), .B(n390), .Y(n613) );
  OR2X1 U640 ( .A(n2394), .B(n391), .Y(n612) );
  OR2X1 U642 ( .A(n2394), .B(n392), .Y(n611) );
  OR2X1 U644 ( .A(n2394), .B(n393), .Y(n610) );
  OR2X1 U646 ( .A(n2394), .B(n394), .Y(n609) );
  OR2X1 U648 ( .A(n2394), .B(n395), .Y(n608) );
  OR2X1 U650 ( .A(n2394), .B(n396), .Y(n607) );
  OR2X1 U652 ( .A(n2394), .B(n397), .Y(n606) );
  OR2X1 U654 ( .A(n2394), .B(n398), .Y(n605) );
  OR2X1 U656 ( .A(n2394), .B(n399), .Y(n604) );
  OR2X1 U658 ( .A(n2394), .B(n400), .Y(n603) );
  OR2X1 U660 ( .A(n2394), .B(n401), .Y(n602) );
  OR2X1 U662 ( .A(n2394), .B(n402), .Y(n601) );
  OR2X1 U664 ( .A(n2394), .B(n403), .Y(n600) );
  OR2X1 U666 ( .A(n2394), .B(n404), .Y(n599) );
  OR2X1 U668 ( .A(n2394), .B(n405), .Y(n598) );
  OR2X1 U670 ( .A(n2394), .B(n406), .Y(n597) );
  OR2X1 U674 ( .A(n2395), .B(n408), .Y(n595) );
  OR2X1 U676 ( .A(n2395), .B(n409), .Y(n594) );
  OR2X1 U678 ( .A(n2395), .B(n410), .Y(n593) );
  OR2X1 U682 ( .A(n2395), .B(n412), .Y(n591) );
  OR2X1 U684 ( .A(n2395), .B(n413), .Y(n590) );
  OR2X1 U686 ( .A(n2395), .B(n414), .Y(n589) );
  OR2X1 U688 ( .A(n2395), .B(n415), .Y(n588) );
  OR2X1 U690 ( .A(n2395), .B(n416), .Y(n587) );
  OR2X1 U692 ( .A(n2395), .B(n417), .Y(n586) );
  OR2X1 U694 ( .A(n2395), .B(n418), .Y(n585) );
  OR2X1 U696 ( .A(n2395), .B(n419), .Y(n584) );
  OR2X1 U698 ( .A(n2395), .B(n420), .Y(n583) );
  OR2X1 U700 ( .A(n2395), .B(n421), .Y(n582) );
  OR2X1 U702 ( .A(n2395), .B(n422), .Y(n581) );
  OR2X1 U704 ( .A(n2395), .B(n423), .Y(n580) );
  OR2X1 U706 ( .A(n2395), .B(n424), .Y(n579) );
  OR2X1 U708 ( .A(n2395), .B(n425), .Y(n578) );
  OR2X1 U710 ( .A(n2395), .B(n426), .Y(n577) );
  OR2X1 U712 ( .A(n2395), .B(n427), .Y(n576) );
  OR2X1 U714 ( .A(n2396), .B(n428), .Y(n575) );
  OR2X1 U716 ( .A(n2396), .B(n429), .Y(n574) );
  OR2X1 U718 ( .A(n2396), .B(n430), .Y(n573) );
  OR2X1 U720 ( .A(n2396), .B(n431), .Y(n572) );
  OR2X1 U722 ( .A(n2396), .B(n432), .Y(n571) );
  OR2X1 U724 ( .A(n2396), .B(n433), .Y(n570) );
  OR2X1 U726 ( .A(n2396), .B(n434), .Y(n569) );
  OR2X1 U730 ( .A(n2396), .B(n436), .Y(n567) );
  OR2X1 U734 ( .A(n2396), .B(n438), .Y(n565) );
  OR2X1 U736 ( .A(n2396), .B(n439), .Y(n564) );
  OR2X1 U738 ( .A(n2396), .B(n440), .Y(n563) );
  OR2X1 U740 ( .A(n2396), .B(n441), .Y(n562) );
  OR2X1 U742 ( .A(n2396), .B(n442), .Y(n561) );
  OR2X1 U744 ( .A(n2396), .B(n443), .Y(n560) );
  OR2X1 U746 ( .A(n2396), .B(n444), .Y(n559) );
  OR2X1 U748 ( .A(n2396), .B(n445), .Y(n558) );
  OR2X1 U750 ( .A(n2396), .B(n446), .Y(n557) );
  OR2X1 U752 ( .A(n2396), .B(n447), .Y(n556) );
  OR2X1 U754 ( .A(n2397), .B(n448), .Y(n555) );
  OR2X1 U758 ( .A(n2397), .B(n450), .Y(n553) );
  OR2X1 U760 ( .A(n2397), .B(n451), .Y(n552) );
  OR2X1 U762 ( .A(n2397), .B(n452), .Y(n551) );
  OR2X1 U776 ( .A(n2397), .B(n459), .Y(n544) );
  OR2X1 U778 ( .A(n2397), .B(n460), .Y(n543) );
  OR2X1 U780 ( .A(n2397), .B(n461), .Y(n542) );
  OR2X1 U782 ( .A(n2397), .B(n462), .Y(n541) );
  OR2X1 U784 ( .A(n2397), .B(n463), .Y(n540) );
  OR2X1 U786 ( .A(n2397), .B(n464), .Y(n539) );
  OR2X1 U790 ( .A(n2397), .B(n466), .Y(n537) );
  OR2X1 U792 ( .A(n2397), .B(n467), .Y(n536) );
  OR2X1 U798 ( .A(n2398), .B(n713), .Y(n533) );
  OR2X1 U800 ( .A(n2398), .B(n712), .Y(n532) );
  OR2X1 U806 ( .A(n2398), .B(n709), .Y(n529) );
  OR2X1 U818 ( .A(n2398), .B(n703), .Y(n523) );
  OR2X1 U820 ( .A(n2398), .B(n702), .Y(n522) );
  OR2X1 U822 ( .A(n2398), .B(n701), .Y(n521) );
  OR2X1 U824 ( .A(n2398), .B(n700), .Y(n520) );
  OR2X1 U828 ( .A(n2398), .B(n698), .Y(n518) );
  OR2X1 U830 ( .A(n2398), .B(n697), .Y(n517) );
  OR2X1 U832 ( .A(n2398), .B(n696), .Y(n516) );
  OR2X1 U834 ( .A(n2399), .B(n695), .Y(n515) );
  OR2X1 U840 ( .A(n2399), .B(n692), .Y(n512) );
  OR2X1 U852 ( .A(n2399), .B(n686), .Y(n506) );
  OR2X1 U856 ( .A(n2399), .B(n684), .Y(n504) );
  OR2X1 U858 ( .A(n2399), .B(n683), .Y(n503) );
  MUX2X1 U862 ( .B(n1057), .A(n1025), .S(n2426), .Y(n861) );
  MUX2X1 U863 ( .B(n1056), .A(n1024), .S(n2426), .Y(n860) );
  MUX2X1 U864 ( .B(n1055), .A(n1023), .S(n2426), .Y(n859) );
  MUX2X1 U865 ( .B(n1054), .A(n1022), .S(n2426), .Y(n858) );
  MUX2X1 U866 ( .B(n1053), .A(n1021), .S(n2426), .Y(n857) );
  MUX2X1 U867 ( .B(n1052), .A(n1020), .S(n2426), .Y(n856) );
  MUX2X1 U868 ( .B(n1051), .A(n1019), .S(n2426), .Y(n855) );
  MUX2X1 U869 ( .B(n1050), .A(n1018), .S(n2426), .Y(n854) );
  MUX2X1 U870 ( .B(n1049), .A(n1017), .S(n2426), .Y(n853) );
  MUX2X1 U871 ( .B(n1048), .A(n1016), .S(n2426), .Y(n852) );
  MUX2X1 U872 ( .B(n1047), .A(n1015), .S(n2426), .Y(n851) );
  MUX2X1 U873 ( .B(n1046), .A(n1014), .S(n2426), .Y(n850) );
  MUX2X1 U874 ( .B(n1045), .A(n1013), .S(n2427), .Y(n849) );
  MUX2X1 U875 ( .B(n1044), .A(n1012), .S(n2427), .Y(n848) );
  MUX2X1 U876 ( .B(n1043), .A(n1011), .S(n2427), .Y(n847) );
  MUX2X1 U877 ( .B(n1042), .A(n1010), .S(n2427), .Y(n846) );
  MUX2X1 U878 ( .B(n1041), .A(n1009), .S(n2427), .Y(n845) );
  MUX2X1 U879 ( .B(n1040), .A(n1008), .S(n2427), .Y(n844) );
  MUX2X1 U880 ( .B(n1039), .A(n1007), .S(n2427), .Y(n843) );
  MUX2X1 U881 ( .B(n1038), .A(n1006), .S(n2427), .Y(n842) );
  MUX2X1 U882 ( .B(n1037), .A(n1005), .S(n2427), .Y(n841) );
  MUX2X1 U883 ( .B(n1036), .A(n1004), .S(n2427), .Y(n840) );
  MUX2X1 U884 ( .B(n1035), .A(n1003), .S(n2427), .Y(n839) );
  MUX2X1 U885 ( .B(n1034), .A(n1002), .S(n2427), .Y(n838) );
  MUX2X1 U886 ( .B(n1033), .A(n1001), .S(n2428), .Y(n837) );
  MUX2X1 U887 ( .B(n1032), .A(n1000), .S(n2428), .Y(n836) );
  MUX2X1 U888 ( .B(n1031), .A(n999), .S(n2428), .Y(n835) );
  MUX2X1 U889 ( .B(n1030), .A(n998), .S(n2428), .Y(n834) );
  MUX2X1 U890 ( .B(n1029), .A(n997), .S(n2428), .Y(n833) );
  MUX2X1 U891 ( .B(n1028), .A(n996), .S(n2428), .Y(n832) );
  MUX2X1 U892 ( .B(n1027), .A(n995), .S(n2428), .Y(n831) );
  MUX2X1 U893 ( .B(n1026), .A(n994), .S(n2428), .Y(n830) );
  MUX2X1 U894 ( .B(n1025), .A(n993), .S(n2428), .Y(n829) );
  MUX2X1 U895 ( .B(n1024), .A(n992), .S(n2428), .Y(n828) );
  MUX2X1 U896 ( .B(n1023), .A(n991), .S(n2428), .Y(n827) );
  MUX2X1 U897 ( .B(n1022), .A(n990), .S(n2428), .Y(n826) );
  MUX2X1 U898 ( .B(n1021), .A(n989), .S(n2429), .Y(n825) );
  MUX2X1 U899 ( .B(n1020), .A(n988), .S(n2429), .Y(n824) );
  MUX2X1 U900 ( .B(n1019), .A(n987), .S(n2429), .Y(n823) );
  MUX2X1 U901 ( .B(n1018), .A(n986), .S(n2429), .Y(n822) );
  MUX2X1 U902 ( .B(n1017), .A(n985), .S(n2429), .Y(n821) );
  MUX2X1 U903 ( .B(n1016), .A(n984), .S(n2429), .Y(n820) );
  MUX2X1 U904 ( .B(n1015), .A(n983), .S(n2429), .Y(n819) );
  MUX2X1 U905 ( .B(n1014), .A(n982), .S(n2429), .Y(n818) );
  MUX2X1 U906 ( .B(n1013), .A(n981), .S(n2429), .Y(n817) );
  MUX2X1 U907 ( .B(n1012), .A(n980), .S(n2429), .Y(n816) );
  MUX2X1 U908 ( .B(n1011), .A(n979), .S(n2429), .Y(n815) );
  MUX2X1 U909 ( .B(n1010), .A(n978), .S(n2429), .Y(n814) );
  MUX2X1 U910 ( .B(n1009), .A(n977), .S(n2430), .Y(n813) );
  MUX2X1 U911 ( .B(n1008), .A(n976), .S(n2430), .Y(n812) );
  MUX2X1 U912 ( .B(n1007), .A(n975), .S(n2430), .Y(n811) );
  MUX2X1 U913 ( .B(n1006), .A(n974), .S(n2430), .Y(n810) );
  MUX2X1 U914 ( .B(n1005), .A(n973), .S(n2430), .Y(n809) );
  MUX2X1 U915 ( .B(n1004), .A(n972), .S(n2430), .Y(n808) );
  MUX2X1 U916 ( .B(n1003), .A(n971), .S(n2430), .Y(n807) );
  MUX2X1 U917 ( .B(n1002), .A(n970), .S(n2430), .Y(n806) );
  MUX2X1 U918 ( .B(n1001), .A(n969), .S(n2430), .Y(n805) );
  MUX2X1 U919 ( .B(n1000), .A(n968), .S(n2430), .Y(n804) );
  MUX2X1 U920 ( .B(n999), .A(n967), .S(n2430), .Y(n803) );
  MUX2X1 U921 ( .B(n998), .A(n966), .S(n2430), .Y(n802) );
  MUX2X1 U922 ( .B(n997), .A(n965), .S(n2336), .Y(n801) );
  MUX2X1 U923 ( .B(n996), .A(n964), .S(n2431), .Y(n800) );
  MUX2X1 U924 ( .B(n995), .A(n963), .S(n2336), .Y(n799) );
  MUX2X1 U925 ( .B(n994), .A(n962), .S(n2433), .Y(n798) );
  MUX2X1 U926 ( .B(n993), .A(n961), .S(n2431), .Y(n797) );
  MUX2X1 U927 ( .B(n992), .A(n960), .S(n2337), .Y(n796) );
  MUX2X1 U928 ( .B(n991), .A(n959), .S(n2432), .Y(n795) );
  MUX2X1 U929 ( .B(n990), .A(n958), .S(n2432), .Y(n794) );
  MUX2X1 U930 ( .B(n989), .A(n957), .S(n2433), .Y(n793) );
  MUX2X1 U931 ( .B(n988), .A(n956), .S(n2431), .Y(n792) );
  MUX2X1 U932 ( .B(n987), .A(n955), .S(n2433), .Y(n791) );
  MUX2X1 U933 ( .B(n986), .A(n954), .S(n2336), .Y(n790) );
  MUX2X1 U934 ( .B(n985), .A(n953), .S(n2337), .Y(n789) );
  MUX2X1 U935 ( .B(n984), .A(n952), .S(n2433), .Y(n788) );
  MUX2X1 U936 ( .B(n983), .A(n951), .S(n2431), .Y(n787) );
  MUX2X1 U937 ( .B(n982), .A(n950), .S(n2336), .Y(n786) );
  MUX2X1 U938 ( .B(n981), .A(n949), .S(n2433), .Y(n785) );
  MUX2X1 U939 ( .B(n980), .A(n948), .S(n2431), .Y(n784) );
  MUX2X1 U940 ( .B(n979), .A(n947), .S(n2433), .Y(n783) );
  MUX2X1 U941 ( .B(n978), .A(n946), .S(n2337), .Y(n782) );
  MUX2X1 U942 ( .B(n977), .A(n945), .S(n2432), .Y(n781) );
  MUX2X1 U943 ( .B(n976), .A(n944), .S(n2432), .Y(n780) );
  MUX2X1 U944 ( .B(n975), .A(n943), .S(n2432), .Y(n779) );
  MUX2X1 U945 ( .B(n974), .A(n942), .S(n2432), .Y(n778) );
  MUX2X1 U946 ( .B(n973), .A(n941), .S(n2336), .Y(n777) );
  MUX2X1 U947 ( .B(n972), .A(n940), .S(n2337), .Y(n776) );
  MUX2X1 U948 ( .B(n971), .A(n939), .S(n2431), .Y(n775) );
  MUX2X1 U949 ( .B(n970), .A(n938), .S(n2336), .Y(n774) );
  MUX2X1 U950 ( .B(n969), .A(n937), .S(n2431), .Y(n773) );
  MUX2X1 U951 ( .B(n968), .A(n936), .S(n2433), .Y(n772) );
  MUX2X1 U952 ( .B(n967), .A(n935), .S(n2431), .Y(n771) );
  MUX2X1 U954 ( .B(n965), .A(n933), .S(n2337), .Y(n769) );
  MUX2X1 U955 ( .B(n964), .A(n932), .S(n2336), .Y(n768) );
  MUX2X1 U956 ( .B(n963), .A(n931), .S(n2337), .Y(n767) );
  MUX2X1 U957 ( .B(n962), .A(n930), .S(n2337), .Y(n766) );
  MUX2X1 U958 ( .B(n961), .A(n929), .S(n2434), .Y(n765) );
  MUX2X1 U959 ( .B(n960), .A(n928), .S(n2434), .Y(n764) );
  MUX2X1 U960 ( .B(n959), .A(n927), .S(n2434), .Y(n763) );
  MUX2X1 U961 ( .B(n958), .A(n926), .S(n2434), .Y(n762) );
  MUX2X1 U962 ( .B(n957), .A(n925), .S(n2434), .Y(n761) );
  MUX2X1 U963 ( .B(n956), .A(n924), .S(n2434), .Y(n760) );
  MUX2X1 U964 ( .B(n955), .A(n923), .S(n2434), .Y(n759) );
  MUX2X1 U965 ( .B(n954), .A(n922), .S(n2434), .Y(n758) );
  MUX2X1 U966 ( .B(n953), .A(n921), .S(n2434), .Y(n757) );
  MUX2X1 U967 ( .B(n952), .A(n920), .S(n2434), .Y(n756) );
  MUX2X1 U968 ( .B(n951), .A(n919), .S(n2434), .Y(n755) );
  MUX2X1 U969 ( .B(n950), .A(n918), .S(n2434), .Y(n754) );
  MUX2X1 U970 ( .B(n949), .A(n917), .S(n2435), .Y(n753) );
  MUX2X1 U971 ( .B(n948), .A(n916), .S(n2435), .Y(n752) );
  MUX2X1 U972 ( .B(n947), .A(n915), .S(n2435), .Y(n751) );
  MUX2X1 U973 ( .B(n946), .A(n914), .S(n2435), .Y(n750) );
  MUX2X1 U974 ( .B(n945), .A(n913), .S(n2435), .Y(n749) );
  MUX2X1 U975 ( .B(n944), .A(n912), .S(n2435), .Y(n748) );
  MUX2X1 U976 ( .B(n943), .A(n911), .S(n2435), .Y(n747) );
  MUX2X1 U977 ( .B(n942), .A(n910), .S(n2435), .Y(n746) );
  MUX2X1 U978 ( .B(n941), .A(n909), .S(n2435), .Y(n745) );
  MUX2X1 U979 ( .B(n940), .A(n2207), .S(n2435), .Y(n744) );
  MUX2X1 U980 ( .B(n939), .A(n907), .S(n2435), .Y(n743) );
  MUX2X1 U981 ( .B(n938), .A(n906), .S(n2435), .Y(n742) );
  MUX2X1 U982 ( .B(n937), .A(n905), .S(n2436), .Y(n741) );
  MUX2X1 U983 ( .B(n936), .A(n904), .S(n2436), .Y(n740) );
  MUX2X1 U984 ( .B(n935), .A(n903), .S(n2436), .Y(n739) );
  MUX2X1 U985 ( .B(n934), .A(n902), .S(n2436), .Y(n738) );
  MUX2X1 U986 ( .B(n933), .A(n901), .S(n2436), .Y(n737) );
  MUX2X1 U987 ( .B(n932), .A(n900), .S(n2436), .Y(n736) );
  MUX2X1 U988 ( .B(n931), .A(n899), .S(n2436), .Y(n735) );
  MUX2X1 U990 ( .B(n929), .A(n897), .S(n2436), .Y(n733) );
  MUX2X1 U991 ( .B(n928), .A(n896), .S(n2436), .Y(n732) );
  MUX2X1 U992 ( .B(n927), .A(n895), .S(n2426), .Y(n731) );
  MUX2X1 U993 ( .B(n926), .A(n894), .S(n2429), .Y(n730) );
  MUX2X1 U994 ( .B(n925), .A(n893), .S(n2437), .Y(n729) );
  MUX2X1 U995 ( .B(n924), .A(n892), .S(n2437), .Y(n728) );
  MUX2X1 U996 ( .B(n923), .A(n891), .S(n2437), .Y(n727) );
  MUX2X1 U997 ( .B(n922), .A(n890), .S(n2437), .Y(n726) );
  MUX2X1 U998 ( .B(n921), .A(n889), .S(n2428), .Y(n725) );
  MUX2X1 U999 ( .B(n920), .A(n888), .S(n2428), .Y(n724) );
  MUX2X1 U1000 ( .B(n919), .A(n887), .S(n2428), .Y(n723) );
  MUX2X1 U1001 ( .B(n918), .A(n886), .S(n2434), .Y(n722) );
  MUX2X1 U1002 ( .B(n917), .A(n885), .S(n2428), .Y(n721) );
  MUX2X1 U1003 ( .B(n916), .A(n884), .S(n2428), .Y(n720) );
  MUX2X1 U1004 ( .B(n915), .A(n883), .S(n2428), .Y(n719) );
  MUX2X1 U1005 ( .B(n914), .A(n882), .S(n2428), .Y(n718) );
  MUX2X1 U1006 ( .B(n913), .A(n881), .S(n2438), .Y(n717) );
  MUX2X1 U1007 ( .B(n912), .A(n880), .S(n2438), .Y(n716) );
  MUX2X1 U1009 ( .B(n910), .A(n878), .S(n2438), .Y(n714) );
  MUX2X1 U1042 ( .B(n1237), .A(n1221), .S(n2448), .Y(n1057) );
  MUX2X1 U1043 ( .B(n1236), .A(n1220), .S(n2448), .Y(n1056) );
  MUX2X1 U1044 ( .B(n1235), .A(n1219), .S(n2448), .Y(n1055) );
  MUX2X1 U1045 ( .B(n1234), .A(n1218), .S(n2448), .Y(n1054) );
  MUX2X1 U1046 ( .B(n1233), .A(n1217), .S(n2448), .Y(n1053) );
  MUX2X1 U1047 ( .B(n1232), .A(n1216), .S(n2448), .Y(n1052) );
  MUX2X1 U1048 ( .B(n1231), .A(n1215), .S(n2448), .Y(n1051) );
  MUX2X1 U1049 ( .B(n1230), .A(n1214), .S(n2448), .Y(n1050) );
  MUX2X1 U1050 ( .B(n1229), .A(n1213), .S(n2448), .Y(n1049) );
  MUX2X1 U1051 ( .B(n1228), .A(n1212), .S(n2448), .Y(n1048) );
  MUX2X1 U1052 ( .B(n1227), .A(n1211), .S(n2448), .Y(n1047) );
  MUX2X1 U1053 ( .B(n1226), .A(n1210), .S(n2448), .Y(n1046) );
  MUX2X1 U1054 ( .B(n1225), .A(n1209), .S(n2449), .Y(n1045) );
  MUX2X1 U1055 ( .B(n1224), .A(n1208), .S(n2449), .Y(n1044) );
  MUX2X1 U1056 ( .B(n1223), .A(n1207), .S(n2449), .Y(n1043) );
  MUX2X1 U1057 ( .B(n1222), .A(n1206), .S(n2449), .Y(n1042) );
  MUX2X1 U1058 ( .B(n1221), .A(n1205), .S(n2449), .Y(n1041) );
  MUX2X1 U1059 ( .B(n1220), .A(n1204), .S(n2449), .Y(n1040) );
  MUX2X1 U1060 ( .B(n1219), .A(n1203), .S(n2449), .Y(n1039) );
  MUX2X1 U1061 ( .B(n1218), .A(n1202), .S(n2449), .Y(n1038) );
  MUX2X1 U1062 ( .B(n1217), .A(n1201), .S(n2449), .Y(n1037) );
  MUX2X1 U1063 ( .B(n1216), .A(n1200), .S(n2449), .Y(n1036) );
  MUX2X1 U1064 ( .B(n1215), .A(n1199), .S(n2449), .Y(n1035) );
  MUX2X1 U1065 ( .B(n1214), .A(n1198), .S(n2449), .Y(n1034) );
  MUX2X1 U1066 ( .B(n1213), .A(n1197), .S(n2450), .Y(n1033) );
  MUX2X1 U1067 ( .B(n1212), .A(n1196), .S(n2450), .Y(n1032) );
  MUX2X1 U1068 ( .B(n1211), .A(n1195), .S(n2450), .Y(n1031) );
  MUX2X1 U1069 ( .B(n1210), .A(n1194), .S(n2450), .Y(n1030) );
  MUX2X1 U1070 ( .B(n1209), .A(n1193), .S(n2450), .Y(n1029) );
  MUX2X1 U1071 ( .B(n1208), .A(n1192), .S(n2450), .Y(n1028) );
  MUX2X1 U1072 ( .B(n1207), .A(n1191), .S(n2450), .Y(n1027) );
  MUX2X1 U1073 ( .B(n1206), .A(n1190), .S(n2450), .Y(n1026) );
  MUX2X1 U1074 ( .B(n1205), .A(n1189), .S(n2450), .Y(n1025) );
  MUX2X1 U1075 ( .B(n1204), .A(n1188), .S(n2450), .Y(n1024) );
  MUX2X1 U1076 ( .B(n1203), .A(n1187), .S(n2450), .Y(n1023) );
  MUX2X1 U1077 ( .B(n1202), .A(n1186), .S(n2450), .Y(n1022) );
  MUX2X1 U1078 ( .B(n1201), .A(n1185), .S(n2451), .Y(n1021) );
  MUX2X1 U1079 ( .B(n1200), .A(n1184), .S(n2451), .Y(n1020) );
  MUX2X1 U1080 ( .B(n1199), .A(n1183), .S(n2451), .Y(n1019) );
  MUX2X1 U1081 ( .B(n1198), .A(n1182), .S(n2451), .Y(n1018) );
  MUX2X1 U1082 ( .B(n1197), .A(n1181), .S(n2451), .Y(n1017) );
  MUX2X1 U1083 ( .B(n1196), .A(n1180), .S(n2451), .Y(n1016) );
  MUX2X1 U1084 ( .B(n1195), .A(n1179), .S(n2451), .Y(n1015) );
  MUX2X1 U1085 ( .B(n1194), .A(n1178), .S(n2451), .Y(n1014) );
  MUX2X1 U1086 ( .B(n1193), .A(n1177), .S(n2451), .Y(n1013) );
  MUX2X1 U1087 ( .B(n1192), .A(n1176), .S(n2451), .Y(n1012) );
  MUX2X1 U1088 ( .B(n1191), .A(n1175), .S(n2451), .Y(n1011) );
  MUX2X1 U1089 ( .B(n1190), .A(n1174), .S(n2451), .Y(n1010) );
  MUX2X1 U1090 ( .B(n1189), .A(n1173), .S(n2452), .Y(n1009) );
  MUX2X1 U1091 ( .B(n1188), .A(n1172), .S(n2452), .Y(n1008) );
  MUX2X1 U1092 ( .B(n1187), .A(n1171), .S(n2452), .Y(n1007) );
  MUX2X1 U1093 ( .B(n1186), .A(n1170), .S(n2452), .Y(n1006) );
  MUX2X1 U1094 ( .B(n1185), .A(n1169), .S(n2452), .Y(n1005) );
  MUX2X1 U1095 ( .B(n1184), .A(n1168), .S(n2452), .Y(n1004) );
  MUX2X1 U1096 ( .B(n1183), .A(n1167), .S(n2452), .Y(n1003) );
  MUX2X1 U1097 ( .B(n1182), .A(n1166), .S(n2452), .Y(n1002) );
  MUX2X1 U1098 ( .B(n1181), .A(n1165), .S(n2452), .Y(n1001) );
  MUX2X1 U1099 ( .B(n1180), .A(n1164), .S(n2452), .Y(n1000) );
  MUX2X1 U1100 ( .B(n1179), .A(n1163), .S(n2452), .Y(n999) );
  MUX2X1 U1101 ( .B(n1178), .A(n1162), .S(n2452), .Y(n998) );
  MUX2X1 U1102 ( .B(n1177), .A(n1161), .S(n2453), .Y(n997) );
  MUX2X1 U1103 ( .B(n1176), .A(n1160), .S(n2453), .Y(n996) );
  MUX2X1 U1104 ( .B(n1175), .A(n1159), .S(n2453), .Y(n995) );
  MUX2X1 U1105 ( .B(n1174), .A(n1158), .S(n2453), .Y(n994) );
  MUX2X1 U1106 ( .B(n1173), .A(n1157), .S(n2453), .Y(n993) );
  MUX2X1 U1107 ( .B(n1172), .A(n1156), .S(n2453), .Y(n992) );
  MUX2X1 U1108 ( .B(n1171), .A(n1155), .S(n2453), .Y(n991) );
  MUX2X1 U1109 ( .B(n1170), .A(n1154), .S(n2453), .Y(n990) );
  MUX2X1 U1110 ( .B(n1169), .A(n1153), .S(n2453), .Y(n989) );
  MUX2X1 U1111 ( .B(n1168), .A(n1152), .S(n2453), .Y(n988) );
  MUX2X1 U1112 ( .B(n1167), .A(n1151), .S(n2453), .Y(n987) );
  MUX2X1 U1113 ( .B(n1166), .A(n1150), .S(n2453), .Y(n986) );
  MUX2X1 U1114 ( .B(n1165), .A(n1149), .S(n2454), .Y(n985) );
  MUX2X1 U1116 ( .B(n1163), .A(n1147), .S(n2456), .Y(n983) );
  MUX2X1 U1117 ( .B(n1162), .A(n1146), .S(n2456), .Y(n982) );
  MUX2X1 U1118 ( .B(n1161), .A(n1145), .S(n2456), .Y(n981) );
  MUX2X1 U1119 ( .B(n1160), .A(n1144), .S(n2455), .Y(n980) );
  MUX2X1 U1120 ( .B(n1159), .A(n1143), .S(n2456), .Y(n979) );
  MUX2X1 U1121 ( .B(n1158), .A(n1142), .S(n2456), .Y(n978) );
  MUX2X1 U1122 ( .B(n1157), .A(n1141), .S(n2454), .Y(n977) );
  MUX2X1 U1124 ( .B(n1155), .A(n1139), .S(n2454), .Y(n975) );
  MUX2X1 U1125 ( .B(n1154), .A(n1138), .S(n2454), .Y(n974) );
  MUX2X1 U1126 ( .B(n1153), .A(n1137), .S(n2455), .Y(n973) );
  MUX2X1 U1127 ( .B(n1152), .A(n1136), .S(n2455), .Y(n972) );
  MUX2X1 U1128 ( .B(n1151), .A(n1135), .S(n2456), .Y(n971) );
  MUX2X1 U1129 ( .B(n1150), .A(n1134), .S(n2456), .Y(n970) );
  MUX2X1 U1130 ( .B(n1149), .A(n1133), .S(n2456), .Y(n969) );
  MUX2X1 U1131 ( .B(n1148), .A(n1132), .S(n2456), .Y(n968) );
  MUX2X1 U1132 ( .B(n1147), .A(n1131), .S(n2455), .Y(n967) );
  MUX2X1 U1133 ( .B(n1146), .A(n1130), .S(n2456), .Y(n966) );
  MUX2X1 U1134 ( .B(n1145), .A(n1129), .S(n2455), .Y(n965) );
  MUX2X1 U1135 ( .B(n1144), .A(n1128), .S(n2456), .Y(n964) );
  MUX2X1 U1136 ( .B(n1143), .A(n1127), .S(n2455), .Y(n963) );
  MUX2X1 U1137 ( .B(n1142), .A(n1126), .S(n2455), .Y(n962) );
  MUX2X1 U1138 ( .B(n1141), .A(n1125), .S(n2455), .Y(n961) );
  MUX2X1 U1139 ( .B(n1140), .A(n1124), .S(n2454), .Y(n960) );
  MUX2X1 U1140 ( .B(n1139), .A(n1123), .S(n2454), .Y(n959) );
  MUX2X1 U1141 ( .B(n1138), .A(n1122), .S(n2454), .Y(n958) );
  MUX2X1 U1142 ( .B(n1137), .A(n1121), .S(n2455), .Y(n957) );
  MUX2X1 U1143 ( .B(n1136), .A(n1120), .S(n2456), .Y(n956) );
  MUX2X1 U1144 ( .B(n1135), .A(n1119), .S(n2455), .Y(n955) );
  MUX2X1 U1145 ( .B(n1134), .A(n1118), .S(n2455), .Y(n954) );
  MUX2X1 U1146 ( .B(n1133), .A(n1117), .S(n2455), .Y(n953) );
  MUX2X1 U1147 ( .B(n1132), .A(n1116), .S(n2456), .Y(n952) );
  MUX2X1 U1148 ( .B(n1131), .A(n1115), .S(n2454), .Y(n951) );
  MUX2X1 U1149 ( .B(n1130), .A(n1114), .S(n2454), .Y(n950) );
  MUX2X1 U1150 ( .B(n1129), .A(n1113), .S(n2457), .Y(n949) );
  MUX2X1 U1151 ( .B(n1128), .A(n1112), .S(n2457), .Y(n948) );
  MUX2X1 U1152 ( .B(n1127), .A(n1111), .S(n2457), .Y(n947) );
  MUX2X1 U1153 ( .B(n1126), .A(n2217), .S(n2457), .Y(n946) );
  MUX2X1 U1154 ( .B(n1125), .A(n1109), .S(n2457), .Y(n945) );
  MUX2X1 U1155 ( .B(n1124), .A(n1108), .S(n2457), .Y(n944) );
  MUX2X1 U1156 ( .B(n1123), .A(n1107), .S(n2457), .Y(n943) );
  MUX2X1 U1158 ( .B(n1121), .A(n1105), .S(n2457), .Y(n941) );
  MUX2X1 U1160 ( .B(n1119), .A(n1103), .S(n2457), .Y(n939) );
  MUX2X1 U1161 ( .B(n1118), .A(n1102), .S(n2457), .Y(n938) );
  MUX2X1 U1162 ( .B(n1117), .A(n1101), .S(n2458), .Y(n937) );
  MUX2X1 U1164 ( .B(n1115), .A(n1099), .S(n2458), .Y(n935) );
  MUX2X1 U1165 ( .B(n1114), .A(n1098), .S(n2458), .Y(n934) );
  MUX2X1 U1166 ( .B(n1113), .A(n1097), .S(n2458), .Y(n933) );
  MUX2X1 U1167 ( .B(n1112), .A(n1096), .S(n2458), .Y(n932) );
  MUX2X1 U1168 ( .B(n1111), .A(n1095), .S(n2458), .Y(n931) );
  MUX2X1 U1169 ( .B(n1110), .A(n1094), .S(n2458), .Y(n930) );
  MUX2X1 U1170 ( .B(n1109), .A(n1093), .S(n2458), .Y(n929) );
  MUX2X1 U1171 ( .B(n1108), .A(n1092), .S(n2458), .Y(n928) );
  MUX2X1 U1172 ( .B(n1107), .A(n1091), .S(n2458), .Y(n927) );
  MUX2X1 U1173 ( .B(n1106), .A(n1090), .S(n2454), .Y(n926) );
  MUX2X1 U1174 ( .B(n1105), .A(n1089), .S(n2459), .Y(n925) );
  MUX2X1 U1175 ( .B(n1104), .A(n2205), .S(n2459), .Y(n924) );
  MUX2X1 U1176 ( .B(n1103), .A(n1087), .S(n2459), .Y(n923) );
  MUX2X1 U1177 ( .B(n1102), .A(n1086), .S(n2459), .Y(n922) );
  MUX2X1 U1178 ( .B(n1101), .A(n1085), .S(n2459), .Y(n921) );
  MUX2X1 U1179 ( .B(n1100), .A(n1084), .S(n2459), .Y(n920) );
  MUX2X1 U1180 ( .B(n1099), .A(n1083), .S(n2459), .Y(n919) );
  MUX2X1 U1181 ( .B(n1098), .A(n1082), .S(n2459), .Y(n918) );
  MUX2X1 U1182 ( .B(n1097), .A(n1081), .S(n2451), .Y(n917) );
  MUX2X1 U1183 ( .B(n1096), .A(n1080), .S(n2459), .Y(n916) );
  MUX2X1 U1184 ( .B(n1095), .A(n1079), .S(n2459), .Y(n915) );
  MUX2X1 U1185 ( .B(n1094), .A(n1078), .S(n2459), .Y(n914) );
  MUX2X1 U1186 ( .B(n1093), .A(n1077), .S(n2460), .Y(n913) );
  MUX2X1 U1187 ( .B(n1092), .A(n1076), .S(n2460), .Y(n912) );
  MUX2X1 U1188 ( .B(n1091), .A(n1075), .S(n2460), .Y(n911) );
  MUX2X1 U1189 ( .B(n1090), .A(n1074), .S(n2460), .Y(n910) );
  MUX2X1 U1190 ( .B(n1089), .A(n1073), .S(n2460), .Y(n909) );
  MUX2X1 U1191 ( .B(n1088), .A(n1072), .S(n2460), .Y(n908) );
  MUX2X1 U1192 ( .B(n1087), .A(n1071), .S(n2460), .Y(n907) );
  MUX2X1 U1193 ( .B(n1086), .A(n1070), .S(n2460), .Y(n906) );
  MUX2X1 U1194 ( .B(n1085), .A(n1069), .S(n2460), .Y(n905) );
  MUX2X1 U1195 ( .B(n1084), .A(n1068), .S(n2460), .Y(n904) );
  MUX2X1 U1196 ( .B(n1083), .A(n1067), .S(n2460), .Y(n903) );
  MUX2X1 U1197 ( .B(n1082), .A(n1066), .S(n2460), .Y(n902) );
  MUX2X1 U1198 ( .B(n1081), .A(n2358), .S(n2461), .Y(n901) );
  MUX2X1 U1202 ( .B(n1077), .A(n2347), .S(n2461), .Y(n897) );
  MUX2X1 U1203 ( .B(n1076), .A(n2350), .S(n2461), .Y(n896) );
  MUX2X1 U1205 ( .B(n1074), .A(n2308), .S(n2461), .Y(n894) );
  MUX2X1 U1238 ( .B(n1421), .A(n1413), .S(n2325), .Y(n1237) );
  MUX2X1 U1239 ( .B(n1420), .A(n1412), .S(n2325), .Y(n1236) );
  MUX2X1 U1240 ( .B(n1419), .A(n1411), .S(n2325), .Y(n1235) );
  MUX2X1 U1241 ( .B(n1418), .A(n1410), .S(n2325), .Y(n1234) );
  MUX2X1 U1242 ( .B(n1417), .A(n1409), .S(n2325), .Y(n1233) );
  MUX2X1 U1243 ( .B(n1416), .A(n1408), .S(n2325), .Y(n1232) );
  MUX2X1 U1244 ( .B(n1415), .A(n1407), .S(n2325), .Y(n1231) );
  MUX2X1 U1245 ( .B(n1414), .A(n1406), .S(n2325), .Y(n1230) );
  MUX2X1 U1246 ( .B(n1413), .A(n1405), .S(n2325), .Y(n1229) );
  MUX2X1 U1247 ( .B(n1412), .A(n1404), .S(n2325), .Y(n1228) );
  MUX2X1 U1248 ( .B(n1411), .A(n1403), .S(n2325), .Y(n1227) );
  MUX2X1 U1249 ( .B(n1410), .A(n1402), .S(n2325), .Y(n1226) );
  MUX2X1 U1250 ( .B(n1409), .A(n1401), .S(n2467), .Y(n1225) );
  MUX2X1 U1251 ( .B(n1408), .A(n1400), .S(n2467), .Y(n1224) );
  MUX2X1 U1252 ( .B(n1407), .A(n1399), .S(n2467), .Y(n1223) );
  MUX2X1 U1253 ( .B(n1406), .A(n1398), .S(n2467), .Y(n1222) );
  MUX2X1 U1254 ( .B(n1405), .A(n1397), .S(n2467), .Y(n1221) );
  MUX2X1 U1255 ( .B(n1404), .A(n1396), .S(n2467), .Y(n1220) );
  MUX2X1 U1256 ( .B(n1403), .A(n1395), .S(n2467), .Y(n1219) );
  MUX2X1 U1257 ( .B(n1402), .A(n1394), .S(n2467), .Y(n1218) );
  MUX2X1 U1258 ( .B(n1401), .A(n1393), .S(n2467), .Y(n1217) );
  MUX2X1 U1259 ( .B(n1400), .A(n1392), .S(n2467), .Y(n1216) );
  MUX2X1 U1260 ( .B(n1399), .A(n1391), .S(n2467), .Y(n1215) );
  MUX2X1 U1261 ( .B(n1398), .A(n1390), .S(n2467), .Y(n1214) );
  MUX2X1 U1262 ( .B(n1397), .A(n1389), .S(n2468), .Y(n1213) );
  MUX2X1 U1263 ( .B(n1396), .A(n1388), .S(n2468), .Y(n1212) );
  MUX2X1 U1264 ( .B(n1395), .A(n1387), .S(n2468), .Y(n1211) );
  MUX2X1 U1265 ( .B(n1394), .A(n1386), .S(n2468), .Y(n1210) );
  MUX2X1 U1266 ( .B(n1393), .A(n1385), .S(n2468), .Y(n1209) );
  MUX2X1 U1267 ( .B(n1392), .A(n1384), .S(n2468), .Y(n1208) );
  MUX2X1 U1268 ( .B(n1391), .A(n1383), .S(n2468), .Y(n1207) );
  MUX2X1 U1269 ( .B(n1390), .A(n1382), .S(n2468), .Y(n1206) );
  MUX2X1 U1270 ( .B(n1389), .A(n1381), .S(n2468), .Y(n1205) );
  MUX2X1 U1271 ( .B(n1388), .A(n1380), .S(n2468), .Y(n1204) );
  MUX2X1 U1272 ( .B(n1387), .A(n1379), .S(n2468), .Y(n1203) );
  MUX2X1 U1273 ( .B(n1386), .A(n1378), .S(n2468), .Y(n1202) );
  MUX2X1 U1274 ( .B(n1385), .A(n1377), .S(n2470), .Y(n1201) );
  MUX2X1 U1275 ( .B(n1384), .A(n1376), .S(n2471), .Y(n1200) );
  MUX2X1 U1276 ( .B(n1383), .A(n1375), .S(n2476), .Y(n1199) );
  MUX2X1 U1277 ( .B(n1382), .A(n1374), .S(n2476), .Y(n1198) );
  MUX2X1 U1278 ( .B(n1381), .A(n1373), .S(n2475), .Y(n1197) );
  MUX2X1 U1279 ( .B(n1380), .A(n1372), .S(n2471), .Y(n1196) );
  MUX2X1 U1280 ( .B(n1379), .A(n1371), .S(n2471), .Y(n1195) );
  MUX2X1 U1281 ( .B(n1378), .A(n1370), .S(n2480), .Y(n1194) );
  MUX2X1 U1282 ( .B(n1377), .A(n1369), .S(n2469), .Y(n1193) );
  MUX2X1 U1283 ( .B(n1376), .A(n1368), .S(n2480), .Y(n1192) );
  MUX2X1 U1284 ( .B(n1375), .A(n1367), .S(n2475), .Y(n1191) );
  MUX2X1 U1285 ( .B(n1374), .A(n1366), .S(n2476), .Y(n1190) );
  MUX2X1 U1286 ( .B(n1373), .A(n1365), .S(n2475), .Y(n1189) );
  MUX2X1 U1287 ( .B(n1372), .A(n1364), .S(n2475), .Y(n1188) );
  MUX2X1 U1288 ( .B(n1371), .A(n1363), .S(n2470), .Y(n1187) );
  MUX2X1 U1289 ( .B(n1370), .A(n1362), .S(n2475), .Y(n1186) );
  MUX2X1 U1290 ( .B(n1369), .A(n1361), .S(n2476), .Y(n1185) );
  MUX2X1 U1291 ( .B(n1368), .A(n1360), .S(n2470), .Y(n1184) );
  MUX2X1 U1292 ( .B(n1367), .A(n1359), .S(n2470), .Y(n1183) );
  MUX2X1 U1293 ( .B(n1366), .A(n1358), .S(n2471), .Y(n1182) );
  MUX2X1 U1294 ( .B(n1365), .A(n1357), .S(n2471), .Y(n1181) );
  MUX2X1 U1295 ( .B(n1364), .A(n1356), .S(n2470), .Y(n1180) );
  MUX2X1 U1296 ( .B(n1363), .A(n1355), .S(n2469), .Y(n1179) );
  MUX2X1 U1297 ( .B(n1362), .A(n1354), .S(n2475), .Y(n1178) );
  MUX2X1 U1298 ( .B(n1361), .A(n1353), .S(n2476), .Y(n1177) );
  MUX2X1 U1299 ( .B(n1360), .A(n1352), .S(n2471), .Y(n1176) );
  MUX2X1 U1300 ( .B(n1359), .A(n1351), .S(n2476), .Y(n1175) );
  MUX2X1 U1301 ( .B(n1358), .A(n1350), .S(n2469), .Y(n1174) );
  MUX2X1 U1302 ( .B(n1357), .A(n1349), .S(n2471), .Y(n1173) );
  MUX2X1 U1303 ( .B(n1356), .A(n1348), .S(n2470), .Y(n1172) );
  MUX2X1 U1304 ( .B(n1355), .A(n1347), .S(n2475), .Y(n1171) );
  MUX2X1 U1305 ( .B(n1354), .A(n1346), .S(n2469), .Y(n1170) );
  MUX2X1 U1306 ( .B(n1353), .A(n1345), .S(n2480), .Y(n1169) );
  MUX2X1 U1307 ( .B(n1352), .A(n1344), .S(n2476), .Y(n1168) );
  MUX2X1 U1308 ( .B(n1351), .A(n1343), .S(n2475), .Y(n1167) );
  MUX2X1 U1309 ( .B(n1350), .A(n1342), .S(n2471), .Y(n1166) );
  MUX2X1 U1310 ( .B(n1349), .A(n1341), .S(n2472), .Y(n1165) );
  MUX2X1 U1311 ( .B(n1348), .A(n1340), .S(n2472), .Y(n1164) );
  MUX2X1 U1312 ( .B(n1347), .A(n1339), .S(n2472), .Y(n1163) );
  MUX2X1 U1313 ( .B(n1346), .A(n1338), .S(n2472), .Y(n1162) );
  MUX2X1 U1314 ( .B(n1345), .A(n1337), .S(n2472), .Y(n1161) );
  MUX2X1 U1315 ( .B(n1344), .A(n1336), .S(n2468), .Y(n1160) );
  MUX2X1 U1316 ( .B(n1343), .A(n1335), .S(n2472), .Y(n1159) );
  MUX2X1 U1317 ( .B(n1342), .A(n1334), .S(n2472), .Y(n1158) );
  MUX2X1 U1318 ( .B(n1341), .A(n1333), .S(n2472), .Y(n1157) );
  MUX2X1 U1319 ( .B(n1340), .A(n1332), .S(n2472), .Y(n1156) );
  MUX2X1 U1320 ( .B(n1339), .A(n1331), .S(n2472), .Y(n1155) );
  MUX2X1 U1321 ( .B(n1338), .A(n1330), .S(n2472), .Y(n1154) );
  MUX2X1 U1322 ( .B(n1337), .A(n1329), .S(n2473), .Y(n1153) );
  MUX2X1 U1323 ( .B(n1336), .A(n1328), .S(n2473), .Y(n1152) );
  MUX2X1 U1324 ( .B(n1335), .A(n1327), .S(n2473), .Y(n1151) );
  MUX2X1 U1325 ( .B(n1334), .A(n1326), .S(n2473), .Y(n1150) );
  MUX2X1 U1326 ( .B(n1333), .A(n1325), .S(n2473), .Y(n1149) );
  MUX2X1 U1327 ( .B(n1332), .A(n1324), .S(n2473), .Y(n1148) );
  MUX2X1 U1328 ( .B(n1331), .A(n1323), .S(n2473), .Y(n1147) );
  MUX2X1 U1329 ( .B(n1330), .A(n1322), .S(n2473), .Y(n1146) );
  MUX2X1 U1330 ( .B(n1329), .A(n1321), .S(n2473), .Y(n1145) );
  MUX2X1 U1331 ( .B(n1328), .A(n1320), .S(n2473), .Y(n1144) );
  MUX2X1 U1332 ( .B(n1327), .A(n1319), .S(n2473), .Y(n1143) );
  MUX2X1 U1333 ( .B(n1326), .A(n1318), .S(n2473), .Y(n1142) );
  MUX2X1 U1334 ( .B(n1325), .A(n1317), .S(n2474), .Y(n1141) );
  MUX2X1 U1335 ( .B(n1324), .A(n1316), .S(n2474), .Y(n1140) );
  MUX2X1 U1336 ( .B(n1323), .A(n1315), .S(n2474), .Y(n1139) );
  MUX2X1 U1337 ( .B(n1322), .A(n1314), .S(n2474), .Y(n1138) );
  MUX2X1 U1338 ( .B(n1321), .A(n1313), .S(n2474), .Y(n1137) );
  MUX2X1 U1339 ( .B(n1320), .A(n1312), .S(n2474), .Y(n1136) );
  MUX2X1 U1340 ( .B(n1319), .A(n1311), .S(n2474), .Y(n1135) );
  MUX2X1 U1341 ( .B(n1318), .A(n1310), .S(n2474), .Y(n1134) );
  MUX2X1 U1342 ( .B(n1317), .A(n1309), .S(n2474), .Y(n1133) );
  MUX2X1 U1343 ( .B(n1316), .A(n1308), .S(n2474), .Y(n1132) );
  MUX2X1 U1344 ( .B(n1315), .A(n1307), .S(n2474), .Y(n1131) );
  MUX2X1 U1345 ( .B(n1314), .A(n1306), .S(n2474), .Y(n1130) );
  MUX2X1 U1346 ( .B(n1313), .A(n1305), .S(n2471), .Y(n1129) );
  MUX2X1 U1347 ( .B(n1312), .A(n1304), .S(n2480), .Y(n1128) );
  MUX2X1 U1348 ( .B(n1311), .A(n1303), .S(n2475), .Y(n1127) );
  MUX2X1 U1349 ( .B(n1310), .A(n1302), .S(n2476), .Y(n1126) );
  MUX2X1 U1350 ( .B(n1309), .A(n1301), .S(n2475), .Y(n1125) );
  MUX2X1 U1351 ( .B(n1308), .A(n1300), .S(n2470), .Y(n1124) );
  MUX2X1 U1352 ( .B(n1307), .A(n1299), .S(n2475), .Y(n1123) );
  MUX2X1 U1353 ( .B(n1306), .A(n1298), .S(n2471), .Y(n1122) );
  MUX2X1 U1354 ( .B(n1305), .A(n1297), .S(n2469), .Y(n1121) );
  MUX2X1 U1355 ( .B(n1304), .A(n1296), .S(n2476), .Y(n1120) );
  MUX2X1 U1356 ( .B(n1303), .A(n1295), .S(n2470), .Y(n1119) );
  MUX2X1 U1357 ( .B(n1302), .A(n1294), .S(n2476), .Y(n1118) );
  MUX2X1 U1358 ( .B(n1301), .A(n1293), .S(n2470), .Y(n1117) );
  MUX2X1 U1359 ( .B(n2330), .A(n1292), .S(n2476), .Y(n1116) );
  MUX2X1 U1360 ( .B(n1299), .A(n1291), .S(n2475), .Y(n1115) );
  MUX2X1 U1361 ( .B(n1298), .A(n1290), .S(n2470), .Y(n1114) );
  MUX2X1 U1362 ( .B(n1297), .A(n1289), .S(n2480), .Y(n1113) );
  MUX2X1 U1363 ( .B(n1296), .A(n1288), .S(n2471), .Y(n1112) );
  MUX2X1 U1364 ( .B(n1295), .A(n1287), .S(n2470), .Y(n1111) );
  MUX2X1 U1365 ( .B(n1294), .A(n1286), .S(n2471), .Y(n1110) );
  MUX2X1 U1366 ( .B(n1293), .A(n1285), .S(n2471), .Y(n1109) );
  MUX2X1 U1367 ( .B(n1292), .A(n1284), .S(n2476), .Y(n1108) );
  MUX2X1 U1368 ( .B(n1291), .A(n1283), .S(n2475), .Y(n1107) );
  MUX2X1 U1369 ( .B(n1290), .A(n1282), .S(n2470), .Y(n1106) );
  MUX2X1 U1370 ( .B(n1289), .A(n1281), .S(n2477), .Y(n1105) );
  MUX2X1 U1371 ( .B(n1288), .A(n1280), .S(n2477), .Y(n1104) );
  MUX2X1 U1372 ( .B(n1287), .A(n1279), .S(n2477), .Y(n1103) );
  MUX2X1 U1373 ( .B(n1286), .A(n1278), .S(n2477), .Y(n1102) );
  MUX2X1 U1374 ( .B(n1285), .A(n1277), .S(n2477), .Y(n1101) );
  MUX2X1 U1375 ( .B(n1284), .A(n1276), .S(n2477), .Y(n1100) );
  MUX2X1 U1376 ( .B(n1283), .A(n1275), .S(n2477), .Y(n1099) );
  MUX2X1 U1377 ( .B(n1282), .A(n1274), .S(n2477), .Y(n1098) );
  MUX2X1 U1378 ( .B(n1281), .A(n1273), .S(n2477), .Y(n1097) );
  MUX2X1 U1379 ( .B(n1280), .A(n1272), .S(n2477), .Y(n1096) );
  MUX2X1 U1380 ( .B(n1279), .A(n1271), .S(n2477), .Y(n1095) );
  MUX2X1 U1381 ( .B(n1278), .A(n1270), .S(n2477), .Y(n1094) );
  MUX2X1 U1382 ( .B(n1277), .A(n1269), .S(n2478), .Y(n1093) );
  MUX2X1 U1383 ( .B(n1276), .A(n1268), .S(n2478), .Y(n1092) );
  MUX2X1 U1384 ( .B(n1275), .A(n1267), .S(n2478), .Y(n1091) );
  MUX2X1 U1385 ( .B(n1274), .A(n1266), .S(n2478), .Y(n1090) );
  MUX2X1 U1386 ( .B(n1273), .A(n1265), .S(n2478), .Y(n1089) );
  MUX2X1 U1388 ( .B(n1271), .A(n1263), .S(n2478), .Y(n1087) );
  MUX2X1 U1389 ( .B(n1270), .A(n1262), .S(n2478), .Y(n1086) );
  MUX2X1 U1390 ( .B(n1269), .A(n1261), .S(n2478), .Y(n1085) );
  MUX2X1 U1391 ( .B(n1268), .A(n1260), .S(n2478), .Y(n1084) );
  MUX2X1 U1392 ( .B(n1267), .A(n1259), .S(n2478), .Y(n1083) );
  MUX2X1 U1393 ( .B(n1266), .A(n1258), .S(n2478), .Y(n1082) );
  MUX2X1 U1394 ( .B(n1265), .A(n1257), .S(n2479), .Y(n1081) );
  MUX2X1 U1395 ( .B(n1264), .A(n1256), .S(n2479), .Y(n1080) );
  MUX2X1 U1396 ( .B(n1263), .A(n1255), .S(n2479), .Y(n1079) );
  MUX2X1 U1397 ( .B(n1262), .A(n1254), .S(n2479), .Y(n1078) );
  MUX2X1 U1398 ( .B(n1261), .A(n1253), .S(n2479), .Y(n1077) );
  MUX2X1 U1399 ( .B(n1260), .A(n1252), .S(n2479), .Y(n1076) );
  MUX2X1 U1400 ( .B(n1259), .A(n1251), .S(n2479), .Y(n1075) );
  MUX2X1 U1401 ( .B(n1258), .A(n1250), .S(n2479), .Y(n1074) );
  MUX2X1 U1402 ( .B(n1257), .A(n1249), .S(n2479), .Y(n1073) );
  MUX2X1 U1403 ( .B(n1256), .A(n1248), .S(n2479), .Y(n1072) );
  MUX2X1 U1404 ( .B(n1255), .A(n1247), .S(n2479), .Y(n1071) );
  MUX2X1 U1406 ( .B(n1253), .A(n1245), .S(n2470), .Y(n1069) );
  MUX2X1 U1407 ( .B(n1252), .A(n1244), .S(n2469), .Y(n1068) );
  MUX2X1 U1408 ( .B(n1251), .A(n1243), .S(n2476), .Y(n1067) );
  MUX2X1 U1409 ( .B(n1250), .A(n1242), .S(n2480), .Y(n1066) );
  MUX2X1 U1418 ( .B(n1601), .A(n1597), .S(n2486), .Y(n1421) );
  MUX2X1 U1419 ( .B(n1600), .A(n1596), .S(n2486), .Y(n1420) );
  MUX2X1 U1420 ( .B(n1599), .A(n1595), .S(n2486), .Y(n1419) );
  MUX2X1 U1421 ( .B(n1598), .A(n1594), .S(n2486), .Y(n1418) );
  MUX2X1 U1422 ( .B(n1597), .A(n1593), .S(n2486), .Y(n1417) );
  MUX2X1 U1423 ( .B(n1596), .A(n1592), .S(n2486), .Y(n1416) );
  MUX2X1 U1424 ( .B(n1595), .A(n1591), .S(n2486), .Y(n1415) );
  MUX2X1 U1425 ( .B(n1594), .A(n1590), .S(n2486), .Y(n1414) );
  MUX2X1 U1426 ( .B(n1593), .A(n1589), .S(n2486), .Y(n1413) );
  MUX2X1 U1427 ( .B(n1592), .A(n1588), .S(n2486), .Y(n1412) );
  MUX2X1 U1428 ( .B(n1591), .A(n1587), .S(n2486), .Y(n1411) );
  MUX2X1 U1429 ( .B(n1590), .A(n1586), .S(n2486), .Y(n1410) );
  MUX2X1 U1430 ( .B(n1589), .A(n1585), .S(n2487), .Y(n1409) );
  MUX2X1 U1431 ( .B(n1588), .A(n1584), .S(n2487), .Y(n1408) );
  MUX2X1 U1432 ( .B(n1587), .A(n1583), .S(n2487), .Y(n1407) );
  MUX2X1 U1433 ( .B(n1586), .A(n1582), .S(n2487), .Y(n1406) );
  MUX2X1 U1434 ( .B(n1585), .A(n1581), .S(n2487), .Y(n1405) );
  MUX2X1 U1435 ( .B(n1584), .A(n1580), .S(n2487), .Y(n1404) );
  MUX2X1 U1436 ( .B(n1583), .A(n1579), .S(n2487), .Y(n1403) );
  MUX2X1 U1437 ( .B(n1582), .A(n1578), .S(n2487), .Y(n1402) );
  MUX2X1 U1438 ( .B(n1581), .A(n1577), .S(n2487), .Y(n1401) );
  MUX2X1 U1439 ( .B(n1580), .A(n1576), .S(n2487), .Y(n1400) );
  MUX2X1 U1440 ( .B(n1579), .A(n1575), .S(n2487), .Y(n1399) );
  MUX2X1 U1441 ( .B(n1578), .A(n1574), .S(n2487), .Y(n1398) );
  MUX2X1 U1442 ( .B(n1577), .A(n1573), .S(n2488), .Y(n1397) );
  MUX2X1 U1443 ( .B(n1576), .A(n1572), .S(n2488), .Y(n1396) );
  MUX2X1 U1444 ( .B(n1575), .A(n1571), .S(n2488), .Y(n1395) );
  MUX2X1 U1445 ( .B(n1574), .A(n1570), .S(n2488), .Y(n1394) );
  MUX2X1 U1446 ( .B(n1573), .A(n1569), .S(n2488), .Y(n1393) );
  MUX2X1 U1447 ( .B(n1572), .A(n1568), .S(n2488), .Y(n1392) );
  MUX2X1 U1448 ( .B(n1571), .A(n1567), .S(n2488), .Y(n1391) );
  MUX2X1 U1449 ( .B(n1570), .A(n1566), .S(n2488), .Y(n1390) );
  MUX2X1 U1450 ( .B(n1569), .A(n1565), .S(n2488), .Y(n1389) );
  MUX2X1 U1451 ( .B(n1568), .A(n1564), .S(n2488), .Y(n1388) );
  MUX2X1 U1452 ( .B(n1567), .A(n1563), .S(n2488), .Y(n1387) );
  MUX2X1 U1453 ( .B(n1566), .A(n1562), .S(n2488), .Y(n1386) );
  MUX2X1 U1454 ( .B(n1565), .A(n1561), .S(n2489), .Y(n1385) );
  MUX2X1 U1455 ( .B(n1564), .A(n1560), .S(n2489), .Y(n1384) );
  MUX2X1 U1456 ( .B(n1563), .A(n1559), .S(n2489), .Y(n1383) );
  MUX2X1 U1457 ( .B(n1562), .A(n1558), .S(n2489), .Y(n1382) );
  MUX2X1 U1458 ( .B(n1561), .A(n1557), .S(n2489), .Y(n1381) );
  MUX2X1 U1459 ( .B(n1560), .A(n1556), .S(n2489), .Y(n1380) );
  MUX2X1 U1460 ( .B(n1559), .A(n1555), .S(n2495), .Y(n1379) );
  MUX2X1 U1461 ( .B(n1558), .A(n1554), .S(n2495), .Y(n1378) );
  MUX2X1 U1462 ( .B(n1557), .A(n1553), .S(n2489), .Y(n1377) );
  MUX2X1 U1463 ( .B(n1556), .A(n1552), .S(n2489), .Y(n1376) );
  MUX2X1 U1464 ( .B(n1555), .A(n1551), .S(n2495), .Y(n1375) );
  MUX2X1 U1465 ( .B(n1554), .A(n1550), .S(n2495), .Y(n1374) );
  MUX2X1 U1466 ( .B(n1553), .A(n1549), .S(n2490), .Y(n1373) );
  MUX2X1 U1467 ( .B(n1552), .A(n1548), .S(n2490), .Y(n1372) );
  MUX2X1 U1468 ( .B(n1551), .A(n1547), .S(n2490), .Y(n1371) );
  MUX2X1 U1469 ( .B(n1550), .A(n1546), .S(n2490), .Y(n1370) );
  MUX2X1 U1470 ( .B(n1549), .A(n1545), .S(n2490), .Y(n1369) );
  MUX2X1 U1471 ( .B(n1548), .A(n1544), .S(n2490), .Y(n1368) );
  MUX2X1 U1472 ( .B(n1547), .A(n1543), .S(n2490), .Y(n1367) );
  MUX2X1 U1473 ( .B(n1546), .A(n1542), .S(n2490), .Y(n1366) );
  MUX2X1 U1474 ( .B(n1545), .A(n1541), .S(n2490), .Y(n1365) );
  MUX2X1 U1475 ( .B(n1544), .A(n1540), .S(n2490), .Y(n1364) );
  MUX2X1 U1476 ( .B(n1543), .A(n1539), .S(n2490), .Y(n1363) );
  MUX2X1 U1477 ( .B(n1542), .A(n1538), .S(n2490), .Y(n1362) );
  MUX2X1 U1478 ( .B(n1541), .A(n1537), .S(n2491), .Y(n1361) );
  MUX2X1 U1479 ( .B(n1540), .A(n1536), .S(n2491), .Y(n1360) );
  MUX2X1 U1480 ( .B(n1539), .A(n1535), .S(n2491), .Y(n1359) );
  MUX2X1 U1481 ( .B(n1538), .A(n1534), .S(n2491), .Y(n1358) );
  MUX2X1 U1482 ( .B(n1537), .A(n1533), .S(n2491), .Y(n1357) );
  MUX2X1 U1483 ( .B(n1536), .A(n1532), .S(n2491), .Y(n1356) );
  MUX2X1 U1484 ( .B(n1535), .A(n1531), .S(n2491), .Y(n1355) );
  MUX2X1 U1485 ( .B(n1534), .A(n1530), .S(n2491), .Y(n1354) );
  MUX2X1 U1486 ( .B(n1533), .A(n1529), .S(n2491), .Y(n1353) );
  MUX2X1 U1487 ( .B(n1532), .A(n1528), .S(n2491), .Y(n1352) );
  MUX2X1 U1488 ( .B(n1531), .A(n1527), .S(n2491), .Y(n1351) );
  MUX2X1 U1489 ( .B(n1530), .A(n1526), .S(n2491), .Y(n1350) );
  MUX2X1 U1490 ( .B(n1529), .A(n1525), .S(n2492), .Y(n1349) );
  MUX2X1 U1491 ( .B(n1528), .A(n1524), .S(n2492), .Y(n1348) );
  MUX2X1 U1492 ( .B(n1527), .A(n1523), .S(n2499), .Y(n1347) );
  MUX2X1 U1493 ( .B(n1526), .A(n1522), .S(n2492), .Y(n1346) );
  MUX2X1 U1494 ( .B(n1525), .A(n1521), .S(n2492), .Y(n1345) );
  MUX2X1 U1495 ( .B(n1524), .A(n1520), .S(n2492), .Y(n1344) );
  MUX2X1 U1496 ( .B(n1523), .A(n1519), .S(n2492), .Y(n1343) );
  MUX2X1 U1497 ( .B(n1522), .A(n1518), .S(n2492), .Y(n1342) );
  MUX2X1 U1498 ( .B(n1521), .A(n1517), .S(n2492), .Y(n1341) );
  MUX2X1 U1499 ( .B(n1520), .A(n1516), .S(n2492), .Y(n1340) );
  MUX2X1 U1500 ( .B(n1519), .A(n1515), .S(n2493), .Y(n1339) );
  MUX2X1 U1501 ( .B(n1518), .A(n1514), .S(n2499), .Y(n1338) );
  MUX2X1 U1502 ( .B(n1517), .A(n1513), .S(n2493), .Y(n1337) );
  MUX2X1 U1503 ( .B(n1516), .A(n1512), .S(n2493), .Y(n1336) );
  MUX2X1 U1504 ( .B(n1515), .A(n1511), .S(n2493), .Y(n1335) );
  MUX2X1 U1505 ( .B(n1514), .A(n1510), .S(n2493), .Y(n1334) );
  MUX2X1 U1506 ( .B(n1513), .A(n1509), .S(n2493), .Y(n1333) );
  MUX2X1 U1507 ( .B(n1512), .A(n1508), .S(n2493), .Y(n1332) );
  MUX2X1 U1508 ( .B(n1511), .A(n1507), .S(n2493), .Y(n1331) );
  MUX2X1 U1509 ( .B(n1510), .A(n1506), .S(n2493), .Y(n1330) );
  MUX2X1 U1510 ( .B(n1509), .A(n1505), .S(n2493), .Y(n1329) );
  MUX2X1 U1511 ( .B(n1508), .A(n1504), .S(n2493), .Y(n1328) );
  MUX2X1 U1512 ( .B(n1507), .A(n1503), .S(n2493), .Y(n1327) );
  MUX2X1 U1513 ( .B(n1506), .A(n1502), .S(n2493), .Y(n1326) );
  MUX2X1 U1514 ( .B(n1505), .A(n1501), .S(n2494), .Y(n1325) );
  MUX2X1 U1515 ( .B(n1504), .A(n1500), .S(n2494), .Y(n1324) );
  MUX2X1 U1516 ( .B(n1503), .A(n1499), .S(n2494), .Y(n1323) );
  MUX2X1 U1517 ( .B(n1502), .A(n1498), .S(n2494), .Y(n1322) );
  MUX2X1 U1518 ( .B(n1501), .A(n1497), .S(n2494), .Y(n1321) );
  MUX2X1 U1519 ( .B(n1500), .A(n1496), .S(n2494), .Y(n1320) );
  MUX2X1 U1520 ( .B(n1499), .A(n1495), .S(n2494), .Y(n1319) );
  MUX2X1 U1521 ( .B(n1498), .A(n1494), .S(n2494), .Y(n1318) );
  MUX2X1 U1522 ( .B(n1497), .A(n1493), .S(n2494), .Y(n1317) );
  MUX2X1 U1523 ( .B(n1496), .A(n1492), .S(n2494), .Y(n1316) );
  MUX2X1 U1524 ( .B(n1495), .A(n1491), .S(n2494), .Y(n1315) );
  MUX2X1 U1525 ( .B(n1494), .A(n1490), .S(n2494), .Y(n1314) );
  MUX2X1 U1526 ( .B(n1493), .A(n1489), .S(n2495), .Y(n1313) );
  MUX2X1 U1527 ( .B(n1492), .A(n1488), .S(n2495), .Y(n1312) );
  MUX2X1 U1528 ( .B(n1491), .A(n1487), .S(n2495), .Y(n1311) );
  MUX2X1 U1529 ( .B(n1490), .A(n1486), .S(n2495), .Y(n1310) );
  MUX2X1 U1530 ( .B(n1489), .A(n1485), .S(n2495), .Y(n1309) );
  MUX2X1 U1531 ( .B(n1488), .A(n1484), .S(n2495), .Y(n1308) );
  MUX2X1 U1532 ( .B(n1487), .A(n1483), .S(n2495), .Y(n1307) );
  MUX2X1 U1533 ( .B(n1486), .A(n1482), .S(n2326), .Y(n1306) );
  MUX2X1 U1534 ( .B(n1485), .A(n1481), .S(n2496), .Y(n1305) );
  MUX2X1 U1535 ( .B(n1484), .A(n1480), .S(n2495), .Y(n1304) );
  MUX2X1 U1536 ( .B(n1483), .A(n1479), .S(n2495), .Y(n1303) );
  MUX2X1 U1537 ( .B(n1482), .A(n1478), .S(n2495), .Y(n1302) );
  MUX2X1 U1538 ( .B(n1481), .A(n1477), .S(n2496), .Y(n1301) );
  MUX2X1 U1539 ( .B(n1480), .A(n1476), .S(n2496), .Y(n1300) );
  MUX2X1 U1540 ( .B(n1479), .A(n1475), .S(n2496), .Y(n1299) );
  MUX2X1 U1541 ( .B(n1478), .A(n1474), .S(n2496), .Y(n1298) );
  MUX2X1 U1542 ( .B(n1477), .A(n1473), .S(n2496), .Y(n1297) );
  MUX2X1 U1543 ( .B(n1476), .A(n1472), .S(n2496), .Y(n1296) );
  MUX2X1 U1544 ( .B(n1475), .A(n1471), .S(n2496), .Y(n1295) );
  MUX2X1 U1545 ( .B(n1474), .A(n1470), .S(n2496), .Y(n1294) );
  MUX2X1 U1546 ( .B(n1473), .A(n1469), .S(n2496), .Y(n1293) );
  MUX2X1 U1547 ( .B(n1472), .A(n1468), .S(n2496), .Y(n1292) );
  MUX2X1 U1548 ( .B(n1471), .A(n1467), .S(n2496), .Y(n1291) );
  MUX2X1 U1549 ( .B(n1470), .A(n1466), .S(n2496), .Y(n1290) );
  MUX2X1 U1550 ( .B(n1469), .A(n1465), .S(n2497), .Y(n1289) );
  MUX2X1 U1551 ( .B(n1468), .A(n1464), .S(n2497), .Y(n1288) );
  MUX2X1 U1552 ( .B(n1467), .A(n1463), .S(n2497), .Y(n1287) );
  MUX2X1 U1553 ( .B(n1466), .A(n1462), .S(n2497), .Y(n1286) );
  MUX2X1 U1554 ( .B(n1465), .A(n1461), .S(n2497), .Y(n1285) );
  MUX2X1 U1555 ( .B(n1464), .A(n1460), .S(n2497), .Y(n1284) );
  MUX2X1 U1556 ( .B(n1463), .A(n1459), .S(n2497), .Y(n1283) );
  MUX2X1 U1557 ( .B(n1462), .A(n1458), .S(n2497), .Y(n1282) );
  MUX2X1 U1558 ( .B(n1461), .A(n1457), .S(n2497), .Y(n1281) );
  MUX2X1 U1559 ( .B(n1460), .A(n1456), .S(n2497), .Y(n1280) );
  MUX2X1 U1560 ( .B(n1459), .A(n1455), .S(n2497), .Y(n1279) );
  MUX2X1 U1561 ( .B(n1458), .A(n1454), .S(n2497), .Y(n1278) );
  MUX2X1 U1562 ( .B(n1457), .A(n1453), .S(n2498), .Y(n1277) );
  MUX2X1 U1563 ( .B(n1456), .A(n1452), .S(n2498), .Y(n1276) );
  MUX2X1 U1564 ( .B(n1455), .A(n1451), .S(n2498), .Y(n1275) );
  MUX2X1 U1565 ( .B(n1454), .A(n1450), .S(n2498), .Y(n1274) );
  MUX2X1 U1566 ( .B(n1453), .A(n1449), .S(n2498), .Y(n1273) );
  MUX2X1 U1567 ( .B(n1452), .A(n1448), .S(n2498), .Y(n1272) );
  MUX2X1 U1568 ( .B(n1451), .A(n1447), .S(n2498), .Y(n1271) );
  MUX2X1 U1569 ( .B(n1450), .A(n1446), .S(n2498), .Y(n1270) );
  MUX2X1 U1570 ( .B(n1449), .A(n1445), .S(n2498), .Y(n1269) );
  MUX2X1 U1571 ( .B(n1448), .A(n1444), .S(n2498), .Y(n1268) );
  MUX2X1 U1572 ( .B(n1447), .A(n1443), .S(n2498), .Y(n1267) );
  MUX2X1 U1573 ( .B(n1446), .A(n1442), .S(n2498), .Y(n1266) );
  MUX2X1 U1574 ( .B(n1445), .A(n1441), .S(n2499), .Y(n1265) );
  MUX2X1 U1575 ( .B(n1444), .A(n1440), .S(n2499), .Y(n1264) );
  MUX2X1 U1578 ( .B(n1441), .A(n1437), .S(n2499), .Y(n1261) );
  MUX2X1 U1580 ( .B(n1439), .A(n1435), .S(n2499), .Y(n1259) );
  MUX2X1 U1581 ( .B(n1438), .A(n1434), .S(n2499), .Y(n1258) );
  MUX2X1 U1582 ( .B(n1437), .A(n1433), .S(n2499), .Y(n1257) );
  MUX2X1 U1583 ( .B(n1436), .A(n1432), .S(n2499), .Y(n1256) );
  MUX2X1 U1584 ( .B(n1435), .A(n1431), .S(n2499), .Y(n1255) );
  MUX2X1 U1585 ( .B(n1434), .A(n1430), .S(n2499), .Y(n1254) );
  MUX2X1 U1586 ( .B(n1433), .A(n1429), .S(n2500), .Y(n1253) );
  MUX2X1 U1587 ( .B(n1432), .A(n1428), .S(n2500), .Y(n1252) );
  MUX2X1 U1588 ( .B(n1431), .A(n1427), .S(n2500), .Y(n1251) );
  MUX2X1 U1589 ( .B(n1430), .A(n1426), .S(n2500), .Y(n1250) );
  MUX2X1 U1590 ( .B(n1429), .A(n1425), .S(n2500), .Y(n1249) );
  MUX2X1 U1591 ( .B(n1428), .A(n1424), .S(n2500), .Y(n1248) );
  MUX2X1 U1592 ( .B(n1427), .A(n2368), .S(n2500), .Y(n1247) );
  MUX2X1 U1593 ( .B(n1426), .A(n2364), .S(n2494), .Y(n1246) );
  MUX2X1 U1602 ( .B(n1781), .A(n1779), .S(n2508), .Y(n1601) );
  MUX2X1 U1603 ( .B(n1780), .A(n1778), .S(n2508), .Y(n1600) );
  MUX2X1 U1604 ( .B(n1779), .A(n1777), .S(n2508), .Y(n1599) );
  MUX2X1 U1605 ( .B(n1778), .A(n1776), .S(n2508), .Y(n1598) );
  MUX2X1 U1606 ( .B(n1777), .A(n1775), .S(n2508), .Y(n1597) );
  MUX2X1 U1607 ( .B(n1776), .A(n1774), .S(n2508), .Y(n1596) );
  MUX2X1 U1608 ( .B(n1775), .A(n1773), .S(n2508), .Y(n1595) );
  MUX2X1 U1609 ( .B(n1774), .A(n1772), .S(n2508), .Y(n1594) );
  MUX2X1 U1610 ( .B(n1773), .A(n1771), .S(n2508), .Y(n1593) );
  MUX2X1 U1611 ( .B(n1772), .A(n1770), .S(n2508), .Y(n1592) );
  MUX2X1 U1612 ( .B(n1771), .A(n1769), .S(n2508), .Y(n1591) );
  MUX2X1 U1613 ( .B(n1770), .A(n1768), .S(n2508), .Y(n1590) );
  MUX2X1 U1614 ( .B(n1769), .A(n1767), .S(n2509), .Y(n1589) );
  MUX2X1 U1615 ( .B(n1768), .A(n1766), .S(n2509), .Y(n1588) );
  MUX2X1 U1616 ( .B(n1767), .A(n1765), .S(n2509), .Y(n1587) );
  MUX2X1 U1617 ( .B(n1766), .A(n1764), .S(n2509), .Y(n1586) );
  MUX2X1 U1618 ( .B(n1765), .A(n1763), .S(n2509), .Y(n1585) );
  MUX2X1 U1619 ( .B(n1764), .A(n1762), .S(n2509), .Y(n1584) );
  MUX2X1 U1620 ( .B(n1763), .A(n1761), .S(n2509), .Y(n1583) );
  MUX2X1 U1621 ( .B(n1762), .A(n1760), .S(n2509), .Y(n1582) );
  MUX2X1 U1622 ( .B(n1761), .A(n1759), .S(n2509), .Y(n1581) );
  MUX2X1 U1623 ( .B(n1760), .A(n1758), .S(n2509), .Y(n1580) );
  MUX2X1 U1624 ( .B(n1759), .A(n1757), .S(n2509), .Y(n1579) );
  MUX2X1 U1625 ( .B(n1758), .A(n1756), .S(n2509), .Y(n1578) );
  MUX2X1 U1626 ( .B(n1757), .A(n1755), .S(n2510), .Y(n1577) );
  MUX2X1 U1627 ( .B(n1756), .A(n1754), .S(n2510), .Y(n1576) );
  MUX2X1 U1628 ( .B(n1755), .A(n1753), .S(n2510), .Y(n1575) );
  MUX2X1 U1629 ( .B(n1754), .A(n1752), .S(n2510), .Y(n1574) );
  MUX2X1 U1630 ( .B(n1753), .A(n1751), .S(n2510), .Y(n1573) );
  MUX2X1 U1631 ( .B(n1752), .A(n1750), .S(n2510), .Y(n1572) );
  MUX2X1 U1632 ( .B(n1751), .A(n1749), .S(n2510), .Y(n1571) );
  MUX2X1 U1633 ( .B(n1750), .A(n1748), .S(n2510), .Y(n1570) );
  MUX2X1 U1634 ( .B(n1749), .A(n1747), .S(n2510), .Y(n1569) );
  MUX2X1 U1635 ( .B(n1748), .A(n1746), .S(n2510), .Y(n1568) );
  MUX2X1 U1636 ( .B(n1747), .A(n1745), .S(n2510), .Y(n1567) );
  MUX2X1 U1637 ( .B(n1746), .A(n1744), .S(n2510), .Y(n1566) );
  MUX2X1 U1638 ( .B(n1745), .A(n1743), .S(n2511), .Y(n1565) );
  MUX2X1 U1639 ( .B(n1744), .A(n1742), .S(n2511), .Y(n1564) );
  MUX2X1 U1640 ( .B(n1743), .A(n1741), .S(n2511), .Y(n1563) );
  MUX2X1 U1641 ( .B(n1742), .A(n1740), .S(n2511), .Y(n1562) );
  MUX2X1 U1642 ( .B(n1741), .A(n1739), .S(n2511), .Y(n1561) );
  MUX2X1 U1643 ( .B(n1740), .A(n1738), .S(n2511), .Y(n1560) );
  MUX2X1 U1644 ( .B(n1739), .A(n1737), .S(n2511), .Y(n1559) );
  MUX2X1 U1645 ( .B(n1738), .A(n1736), .S(n2511), .Y(n1558) );
  MUX2X1 U1646 ( .B(n1737), .A(n1735), .S(n2511), .Y(n1557) );
  MUX2X1 U1647 ( .B(n1736), .A(n1734), .S(n2511), .Y(n1556) );
  MUX2X1 U1648 ( .B(n1735), .A(n1733), .S(n2511), .Y(n1555) );
  MUX2X1 U1649 ( .B(n1734), .A(n1732), .S(n2511), .Y(n1554) );
  MUX2X1 U1650 ( .B(n1733), .A(n1731), .S(n2512), .Y(n1553) );
  MUX2X1 U1651 ( .B(n1732), .A(n1730), .S(n2512), .Y(n1552) );
  MUX2X1 U1652 ( .B(n1731), .A(n1729), .S(n2512), .Y(n1551) );
  MUX2X1 U1653 ( .B(n1730), .A(n1728), .S(n2512), .Y(n1550) );
  MUX2X1 U1654 ( .B(n1729), .A(n1727), .S(n2512), .Y(n1549) );
  MUX2X1 U1655 ( .B(n1728), .A(n1726), .S(n2512), .Y(n1548) );
  MUX2X1 U1656 ( .B(n1727), .A(n1725), .S(n2512), .Y(n1547) );
  MUX2X1 U1657 ( .B(n1726), .A(n1724), .S(n2512), .Y(n1546) );
  MUX2X1 U1658 ( .B(n1725), .A(n1723), .S(n2512), .Y(n1545) );
  MUX2X1 U1659 ( .B(n1724), .A(n1722), .S(n2512), .Y(n1544) );
  MUX2X1 U1660 ( .B(n1723), .A(n1721), .S(n2512), .Y(n1543) );
  MUX2X1 U1661 ( .B(n1722), .A(n1720), .S(n2512), .Y(n1542) );
  MUX2X1 U1662 ( .B(n1721), .A(n1719), .S(n2513), .Y(n1541) );
  MUX2X1 U1663 ( .B(n1720), .A(n1718), .S(n2513), .Y(n1540) );
  MUX2X1 U1664 ( .B(n1719), .A(n1717), .S(n2513), .Y(n1539) );
  MUX2X1 U1665 ( .B(n1718), .A(n1716), .S(n2513), .Y(n1538) );
  MUX2X1 U1666 ( .B(n1717), .A(n1715), .S(n2513), .Y(n1537) );
  MUX2X1 U1667 ( .B(n1716), .A(n1714), .S(n2513), .Y(n1536) );
  MUX2X1 U1668 ( .B(n1715), .A(n1713), .S(n2513), .Y(n1535) );
  MUX2X1 U1669 ( .B(n1714), .A(n1712), .S(n2513), .Y(n1534) );
  MUX2X1 U1670 ( .B(n1713), .A(n1711), .S(n2513), .Y(n1533) );
  MUX2X1 U1671 ( .B(n1712), .A(n1710), .S(n2513), .Y(n1532) );
  MUX2X1 U1672 ( .B(n1711), .A(n1709), .S(n2513), .Y(n1531) );
  MUX2X1 U1673 ( .B(n1710), .A(n1708), .S(n2513), .Y(n1530) );
  MUX2X1 U1674 ( .B(n1709), .A(n1707), .S(n2514), .Y(n1529) );
  MUX2X1 U1675 ( .B(n1708), .A(n1706), .S(n2514), .Y(n1528) );
  MUX2X1 U1676 ( .B(n1707), .A(n1705), .S(n2514), .Y(n1527) );
  MUX2X1 U1677 ( .B(n1706), .A(n1704), .S(n2514), .Y(n1526) );
  MUX2X1 U1678 ( .B(n1705), .A(n1703), .S(n2514), .Y(n1525) );
  MUX2X1 U1679 ( .B(n1704), .A(n1702), .S(n2514), .Y(n1524) );
  MUX2X1 U1680 ( .B(n1703), .A(n1701), .S(n2514), .Y(n1523) );
  MUX2X1 U1682 ( .B(n1701), .A(n1699), .S(n2514), .Y(n1521) );
  MUX2X1 U1683 ( .B(n1700), .A(n1698), .S(n2514), .Y(n1520) );
  MUX2X1 U1684 ( .B(n1699), .A(n1697), .S(n2514), .Y(n1519) );
  MUX2X1 U1685 ( .B(n1698), .A(n1696), .S(n2514), .Y(n1518) );
  MUX2X1 U1686 ( .B(n1697), .A(n1695), .S(n2515), .Y(n1517) );
  MUX2X1 U1687 ( .B(n1696), .A(n1694), .S(n2515), .Y(n1516) );
  MUX2X1 U1688 ( .B(n1695), .A(n1693), .S(n2515), .Y(n1515) );
  MUX2X1 U1689 ( .B(n1694), .A(n1692), .S(n2515), .Y(n1514) );
  MUX2X1 U1690 ( .B(n1693), .A(n1691), .S(n2515), .Y(n1513) );
  MUX2X1 U1691 ( .B(n1692), .A(n1690), .S(n2515), .Y(n1512) );
  MUX2X1 U1692 ( .B(n1691), .A(n1689), .S(n2515), .Y(n1511) );
  MUX2X1 U1693 ( .B(n1690), .A(n1688), .S(n2515), .Y(n1510) );
  MUX2X1 U1694 ( .B(n1689), .A(n1687), .S(n2515), .Y(n1509) );
  MUX2X1 U1695 ( .B(n1688), .A(n1686), .S(n2515), .Y(n1508) );
  MUX2X1 U1696 ( .B(n1687), .A(n1685), .S(n2515), .Y(n1507) );
  MUX2X1 U1697 ( .B(n1686), .A(n1684), .S(n2515), .Y(n1506) );
  MUX2X1 U1698 ( .B(n1685), .A(n1683), .S(n2321), .Y(n1505) );
  MUX2X1 U1699 ( .B(n1684), .A(n1682), .S(n2321), .Y(n1504) );
  MUX2X1 U1700 ( .B(n1683), .A(n1681), .S(n2321), .Y(n1503) );
  MUX2X1 U1701 ( .B(n1682), .A(n1680), .S(n2321), .Y(n1502) );
  MUX2X1 U1702 ( .B(n1681), .A(n1679), .S(n2516), .Y(n1501) );
  MUX2X1 U1703 ( .B(n1680), .A(n1678), .S(n2321), .Y(n1500) );
  MUX2X1 U1704 ( .B(n1679), .A(n1677), .S(n2516), .Y(n1499) );
  MUX2X1 U1705 ( .B(n1678), .A(n1676), .S(n2516), .Y(n1498) );
  MUX2X1 U1706 ( .B(n1677), .A(n1675), .S(n2516), .Y(n1497) );
  MUX2X1 U1707 ( .B(n1676), .A(n1674), .S(n2516), .Y(n1496) );
  MUX2X1 U1708 ( .B(n1675), .A(n1673), .S(n2516), .Y(n1495) );
  MUX2X1 U1709 ( .B(n1674), .A(n1672), .S(n2321), .Y(n1494) );
  MUX2X1 U1710 ( .B(n1673), .A(n1671), .S(n2517), .Y(n1493) );
  MUX2X1 U1711 ( .B(n1672), .A(n1670), .S(n2517), .Y(n1492) );
  MUX2X1 U1712 ( .B(n1671), .A(n1669), .S(n2517), .Y(n1491) );
  MUX2X1 U1713 ( .B(n1670), .A(n1668), .S(n2517), .Y(n1490) );
  MUX2X1 U1714 ( .B(n1669), .A(n1667), .S(n2517), .Y(n1489) );
  MUX2X1 U1715 ( .B(n1668), .A(n1666), .S(n2517), .Y(n1488) );
  MUX2X1 U1716 ( .B(n1667), .A(n1665), .S(n2517), .Y(n1487) );
  MUX2X1 U1717 ( .B(n1666), .A(n1664), .S(n2517), .Y(n1486) );
  MUX2X1 U1718 ( .B(n1665), .A(n1663), .S(n2517), .Y(n1485) );
  MUX2X1 U1719 ( .B(n1664), .A(n1662), .S(n2517), .Y(n1484) );
  MUX2X1 U1720 ( .B(n1663), .A(n1661), .S(n2517), .Y(n1483) );
  MUX2X1 U1721 ( .B(n1662), .A(n1660), .S(n2520), .Y(n1482) );
  MUX2X1 U1722 ( .B(n1661), .A(n1659), .S(n2518), .Y(n1481) );
  MUX2X1 U1723 ( .B(n1660), .A(n1658), .S(n2518), .Y(n1480) );
  MUX2X1 U1724 ( .B(n1659), .A(n1657), .S(n2518), .Y(n1479) );
  MUX2X1 U1725 ( .B(n1658), .A(n1656), .S(n2518), .Y(n1478) );
  MUX2X1 U1726 ( .B(n1657), .A(n1655), .S(n2518), .Y(n1477) );
  MUX2X1 U1728 ( .B(n1655), .A(n1653), .S(n2518), .Y(n1475) );
  MUX2X1 U1730 ( .B(n1653), .A(n1651), .S(n2518), .Y(n1473) );
  MUX2X1 U1731 ( .B(n1652), .A(n1650), .S(n2518), .Y(n1472) );
  MUX2X1 U1732 ( .B(n1651), .A(n1649), .S(n2518), .Y(n1471) );
  MUX2X1 U1733 ( .B(n1650), .A(n1648), .S(n2518), .Y(n1470) );
  MUX2X1 U1734 ( .B(n1649), .A(n1647), .S(n2519), .Y(n1469) );
  MUX2X1 U1735 ( .B(n1648), .A(n1646), .S(n2519), .Y(n1468) );
  MUX2X1 U1736 ( .B(n1647), .A(n1645), .S(n2519), .Y(n1467) );
  MUX2X1 U1738 ( .B(n1645), .A(n1643), .S(n2519), .Y(n1465) );
  MUX2X1 U1739 ( .B(n1644), .A(n1642), .S(n2519), .Y(n1464) );
  MUX2X1 U1740 ( .B(n1643), .A(n1641), .S(n2519), .Y(n1463) );
  MUX2X1 U1741 ( .B(n1642), .A(n1640), .S(n2519), .Y(n1462) );
  MUX2X1 U1742 ( .B(n1641), .A(n1639), .S(n2519), .Y(n1461) );
  MUX2X1 U1743 ( .B(n1640), .A(n1638), .S(n2519), .Y(n1460) );
  MUX2X1 U1744 ( .B(n1639), .A(n1637), .S(n2519), .Y(n1459) );
  MUX2X1 U1745 ( .B(n1638), .A(n1636), .S(n2519), .Y(n1458) );
  MUX2X1 U1746 ( .B(n1637), .A(n1635), .S(n2520), .Y(n1457) );
  MUX2X1 U1747 ( .B(n1636), .A(n1634), .S(n2520), .Y(n1456) );
  MUX2X1 U1748 ( .B(n1635), .A(n1633), .S(n2520), .Y(n1455) );
  MUX2X1 U1749 ( .B(n1634), .A(n1632), .S(n2520), .Y(n1454) );
  MUX2X1 U1750 ( .B(n1633), .A(n1631), .S(n2520), .Y(n1453) );
  MUX2X1 U1751 ( .B(n1632), .A(n1630), .S(n2520), .Y(n1452) );
  MUX2X1 U1752 ( .B(n1631), .A(n1629), .S(n2520), .Y(n1451) );
  MUX2X1 U1753 ( .B(n1630), .A(n1628), .S(n2520), .Y(n1450) );
  MUX2X1 U1754 ( .B(n1629), .A(n1627), .S(n2520), .Y(n1449) );
  MUX2X1 U1755 ( .B(n1628), .A(n1626), .S(n2520), .Y(n1448) );
  MUX2X1 U1756 ( .B(n1627), .A(n1625), .S(n2520), .Y(n1447) );
  MUX2X1 U1757 ( .B(n1626), .A(n1624), .S(n2520), .Y(n1446) );
  MUX2X1 U1758 ( .B(n1625), .A(n1623), .S(n2521), .Y(n1445) );
  MUX2X1 U1759 ( .B(n1624), .A(n1622), .S(n2521), .Y(n1444) );
  MUX2X1 U1760 ( .B(n1623), .A(n1621), .S(n2521), .Y(n1443) );
  MUX2X1 U1762 ( .B(n1621), .A(n1619), .S(n2521), .Y(n1441) );
  MUX2X1 U1763 ( .B(n1620), .A(n1618), .S(n2521), .Y(n1440) );
  MUX2X1 U1764 ( .B(n1619), .A(n1617), .S(n2521), .Y(n1439) );
  MUX2X1 U1765 ( .B(n1618), .A(n1616), .S(n2521), .Y(n1438) );
  MUX2X1 U1766 ( .B(n1617), .A(n1615), .S(n2521), .Y(n1437) );
  MUX2X1 U1767 ( .B(n1616), .A(n1614), .S(n2521), .Y(n1436) );
  MUX2X1 U1768 ( .B(n1615), .A(n1613), .S(n2521), .Y(n1435) );
  MUX2X1 U1770 ( .B(n1613), .A(n1611), .S(n2522), .Y(n1433) );
  MUX2X1 U1771 ( .B(n1612), .A(n1610), .S(n2522), .Y(n1432) );
  MUX2X1 U1772 ( .B(n1611), .A(n1609), .S(n2522), .Y(n1431) );
  MUX2X1 U1773 ( .B(n1610), .A(n1608), .S(n2522), .Y(n1430) );
  MUX2X1 U1774 ( .B(n1609), .A(n1607), .S(n2522), .Y(n1429) );
  MUX2X1 U1776 ( .B(n1607), .A(n1605), .S(n2522), .Y(n1427) );
  MUX2X1 U1777 ( .B(n1606), .A(n1604), .S(n2522), .Y(n1426) );
  MUX2X1 U1778 ( .B(n1605), .A(n1603), .S(n2522), .Y(n1425) );
  MUX2X1 U1779 ( .B(n1604), .A(n1602), .S(n2522), .Y(n1424) );
  MUX2X1 U1988 ( .B(n1606), .A(n1608), .S(n2523), .Y(n1428) );
  MUX2X1 U1989 ( .B(n1080), .A(n2361), .S(n2202), .Y(n900) );
  INVX8 U1990 ( .A(n2334), .Y(n2202) );
  INVX4 U1991 ( .A(n2523), .Y(n2522) );
  OR2X2 U1992 ( .A(n2398), .B(n710), .Y(n530) );
  OR2X1 U1993 ( .A(n2399), .B(n2418), .Y(n2203) );
  INVX4 U1994 ( .A(n2419), .Y(n2418) );
  AND2X2 U1995 ( .A(n2262), .B(n2229), .Y(n2378) );
  INVX1 U1996 ( .A(n2386), .Y(n2225) );
  INVX4 U1997 ( .A(n2222), .Y(n2380) );
  OR2X2 U1998 ( .A(SH[21]), .B(SH[26]), .Y(n2323) );
  INVX4 U1999 ( .A(n2386), .Y(n2315) );
  INVX2 U2000 ( .A(n2294), .Y(n2316) );
  OR2X1 U2001 ( .A(SH[31]), .B(SH[17]), .Y(n2319) );
  OR2X1 U2002 ( .A(SH[19]), .B(SH[18]), .Y(n2376) );
  INVX1 U2003 ( .A(n2214), .Y(n899) );
  INVX1 U2004 ( .A(n1079), .Y(n2215) );
  INVX1 U2005 ( .A(n723), .Y(n460) );
  INVX1 U2006 ( .A(n2210), .Y(n554) );
  INVX1 U2007 ( .A(n1075), .Y(n2213) );
  INVX1 U2008 ( .A(n714), .Y(n469) );
  INVX1 U2009 ( .A(n2442), .Y(n2432) );
  INVX1 U2010 ( .A(n722), .Y(n461) );
  INVX1 U2011 ( .A(n1088), .Y(n2204) );
  INVX1 U2012 ( .A(n2204), .Y(n2205) );
  INVX1 U2013 ( .A(n908), .Y(n2206) );
  INVX1 U2014 ( .A(n2206), .Y(n2207) );
  OR2X2 U2015 ( .A(n2399), .B(n694), .Y(n514) );
  OR2X2 U2016 ( .A(n514), .B(n2418), .Y(n206) );
  OR2X2 U2017 ( .A(n2398), .B(n705), .Y(n525) );
  OR2X2 U2018 ( .A(n2398), .B(n706), .Y(n526) );
  MUX2X1 U2019 ( .B(n1439), .A(n1443), .S(n2501), .Y(n1263) );
  INVX8 U2020 ( .A(n2501), .Y(n2499) );
  OR2X1 U2021 ( .A(n2480), .B(n2462), .Y(n2208) );
  OR2X2 U2022 ( .A(n2500), .B(n1239), .Y(n1244) );
  OR2X2 U2023 ( .A(n2398), .B(n704), .Y(n524) );
  OR2X2 U2024 ( .A(n524), .B(n2417), .Y(n216) );
  MUX2X1 U2025 ( .B(n879), .A(n911), .S(n2440), .Y(n715) );
  INVX8 U2026 ( .A(n2440), .Y(n2438) );
  OR2X1 U2027 ( .A(n2397), .B(n2416), .Y(n2209) );
  AND2X2 U2028 ( .A(n2402), .B(n734), .Y(n2210) );
  MUX2X1 U2029 ( .B(n1426), .A(n2364), .S(n2494), .Y(n2211) );
  MUX2X1 U2030 ( .B(n2211), .A(n1254), .S(n2481), .Y(n1070) );
  INVX2 U2031 ( .A(n1422), .Y(n2364) );
  INVX8 U2032 ( .A(n2481), .Y(n2479) );
  MUX2X1 U2033 ( .B(n930), .A(n898), .S(n2432), .Y(n734) );
  INVX1 U2034 ( .A(n1078), .Y(n2220) );
  INVX1 U2035 ( .A(n2219), .Y(n898) );
  MUX2X1 U2036 ( .B(n1059), .A(n2213), .S(n2463), .Y(n2212) );
  INVX1 U2037 ( .A(n2212), .Y(n895) );
  INVX4 U2038 ( .A(n2463), .Y(n2461) );
  OR2X2 U2039 ( .A(n2399), .B(n685), .Y(n505) );
  OR2X2 U2040 ( .A(n2203), .B(n685), .Y(n197) );
  OR2X2 U2041 ( .A(n2398), .B(n707), .Y(n527) );
  OR2X2 U2042 ( .A(n2398), .B(n468), .Y(n535) );
  MUX2X1 U2043 ( .B(n2215), .A(n1063), .S(n2461), .Y(n2214) );
  MUX2X1 U2044 ( .B(n1652), .A(n1654), .S(n2507), .Y(n1474) );
  INVX1 U2045 ( .A(n1110), .Y(n2216) );
  INVX1 U2046 ( .A(n2216), .Y(n2217) );
  INVX1 U2047 ( .A(n715), .Y(n468) );
  AND2X2 U2048 ( .A(n349), .B(n2384), .Y(B[155]) );
  OR2X2 U2049 ( .A(n2500), .B(n1238), .Y(n1245) );
  OR2X2 U2050 ( .A(n2500), .B(n2476), .Y(n2218) );
  INVX4 U2051 ( .A(n2224), .Y(n2333) );
  OR2X1 U2052 ( .A(n550), .B(n2416), .Y(n242) );
  MUX2X1 U2053 ( .B(n1062), .A(n2220), .S(n2463), .Y(n2219) );
  INVX2 U2054 ( .A(n2441), .Y(n2436) );
  INVX1 U2055 ( .A(n2385), .Y(n2221) );
  INVX1 U2056 ( .A(n1782), .Y(n2222) );
  INVX2 U2057 ( .A(n2385), .Y(n2223) );
  INVX1 U2058 ( .A(n1782), .Y(n2224) );
  OR2X2 U2059 ( .A(n2397), .B(n453), .Y(n550) );
  AND2X2 U2060 ( .A(n347), .B(n2316), .Y(B[153]) );
  AND2X2 U2061 ( .A(n353), .B(n2316), .Y(B[159]) );
  INVX8 U2062 ( .A(n2293), .Y(n2381) );
  OR2X2 U2063 ( .A(SH[23]), .B(SH[22]), .Y(n1794) );
  OR2X2 U2064 ( .A(SH[16]), .B(SH[10]), .Y(n1803) );
  AND2X2 U2065 ( .A(n343), .B(n2316), .Y(B[149]) );
  AND2X2 U2066 ( .A(n299), .B(n2379), .Y(B[105]) );
  AND2X2 U2067 ( .A(n2327), .B(n1784), .Y(n2226) );
  AND2X2 U2068 ( .A(n268), .B(n2384), .Y(B[74]) );
  INVX1 U2069 ( .A(n2385), .Y(n2331) );
  INVX1 U2070 ( .A(n2335), .Y(n2227) );
  OR2X1 U2071 ( .A(n2209), .B(n449), .Y(n246) );
  INVX1 U2072 ( .A(n246), .Y(n2228) );
  OR2X2 U2073 ( .A(n1804), .B(SH[11]), .Y(n2320) );
  INVX1 U2074 ( .A(n2320), .Y(n2229) );
  OR2X2 U2075 ( .A(n1422), .B(n2218), .Y(n2322) );
  AND2X2 U2076 ( .A(n1784), .B(n2327), .Y(n1782) );
  OR2X2 U2077 ( .A(n879), .B(n2439), .Y(n683) );
  OR2X2 U2078 ( .A(n880), .B(n2439), .Y(n684) );
  OR2X2 U2079 ( .A(n881), .B(n2439), .Y(n685) );
  OR2X2 U2080 ( .A(n889), .B(n2439), .Y(n693) );
  OR2X1 U2081 ( .A(n897), .B(n2438), .Y(n701) );
  INVX1 U2082 ( .A(n701), .Y(n2230) );
  OR2X2 U2083 ( .A(n905), .B(n2438), .Y(n709) );
  OR2X1 U2084 ( .A(n503), .B(n2418), .Y(n195) );
  INVX1 U2085 ( .A(n195), .Y(n2231) );
  OR2X2 U2086 ( .A(n504), .B(n2418), .Y(n196) );
  INVX1 U2087 ( .A(n196), .Y(n2232) );
  INVX1 U2088 ( .A(n197), .Y(n2233) );
  OR2X1 U2089 ( .A(n511), .B(n2418), .Y(n203) );
  INVX1 U2090 ( .A(n203), .Y(n2234) );
  OR2X1 U2091 ( .A(n512), .B(n2418), .Y(n204) );
  INVX1 U2092 ( .A(n204), .Y(n2235) );
  INVX1 U2093 ( .A(n206), .Y(n2236) );
  OR2X1 U2094 ( .A(n518), .B(n2417), .Y(n210) );
  INVX1 U2095 ( .A(n210), .Y(n2237) );
  OR2X2 U2096 ( .A(n526), .B(n2417), .Y(n218) );
  INVX1 U2097 ( .A(n218), .Y(n2238) );
  OR2X2 U2098 ( .A(n527), .B(n2417), .Y(n219) );
  INVX1 U2099 ( .A(n219), .Y(n2239) );
  OR2X2 U2100 ( .A(n528), .B(n2417), .Y(n220) );
  INVX1 U2101 ( .A(n220), .Y(n2240) );
  OR2X2 U2102 ( .A(n529), .B(n2417), .Y(n221) );
  INVX1 U2103 ( .A(n221), .Y(n2241) );
  OR2X1 U2104 ( .A(n532), .B(n2417), .Y(n224) );
  INVX1 U2105 ( .A(n224), .Y(n2242) );
  OR2X2 U2106 ( .A(n536), .B(n2417), .Y(n228) );
  INVX1 U2107 ( .A(n228), .Y(n2243) );
  OR2X1 U2108 ( .A(n537), .B(n2417), .Y(n229) );
  INVX1 U2109 ( .A(n229), .Y(n2244) );
  OR2X1 U2110 ( .A(n539), .B(n2416), .Y(n231) );
  INVX1 U2111 ( .A(n231), .Y(n2245) );
  OR2X1 U2112 ( .A(n540), .B(n2416), .Y(n232) );
  INVX1 U2113 ( .A(n232), .Y(n2246) );
  OR2X1 U2114 ( .A(n541), .B(n2416), .Y(n233) );
  INVX1 U2115 ( .A(n233), .Y(n2247) );
  OR2X1 U2116 ( .A(n542), .B(n2416), .Y(n234) );
  INVX1 U2117 ( .A(n234), .Y(n2248) );
  OR2X1 U2118 ( .A(n543), .B(n2416), .Y(n235) );
  INVX1 U2119 ( .A(n235), .Y(n2249) );
  OR2X1 U2120 ( .A(n544), .B(n2416), .Y(n236) );
  INVX1 U2121 ( .A(n236), .Y(n2250) );
  OR2X1 U2122 ( .A(n545), .B(n2416), .Y(n237) );
  INVX1 U2123 ( .A(n237), .Y(n2251) );
  INVX1 U2124 ( .A(n242), .Y(n2252) );
  OR2X2 U2125 ( .A(n552), .B(n2416), .Y(n244) );
  INVX1 U2126 ( .A(n244), .Y(n2253) );
  OR2X1 U2127 ( .A(n555), .B(n2416), .Y(n247) );
  INVX1 U2128 ( .A(n247), .Y(n2254) );
  OR2X2 U2129 ( .A(n557), .B(n2416), .Y(n249) );
  INVX1 U2130 ( .A(n249), .Y(n2255) );
  OR2X2 U2131 ( .A(n558), .B(n2416), .Y(n250) );
  INVX1 U2132 ( .A(n250), .Y(n2256) );
  OR2X1 U2133 ( .A(n559), .B(n2415), .Y(n251) );
  INVX1 U2134 ( .A(n251), .Y(n2257) );
  OR2X1 U2135 ( .A(n560), .B(n2415), .Y(n252) );
  INVX1 U2136 ( .A(n252), .Y(n2258) );
  OR2X1 U2137 ( .A(n561), .B(n2415), .Y(n253) );
  INVX1 U2138 ( .A(n253), .Y(n2259) );
  OR2X2 U2139 ( .A(n562), .B(n2415), .Y(n254) );
  INVX1 U2140 ( .A(n254), .Y(n2260) );
  OR2X1 U2141 ( .A(n563), .B(n2415), .Y(n255) );
  INVX1 U2142 ( .A(n255), .Y(n2261) );
  INVX1 U2143 ( .A(n2319), .Y(n2262) );
  INVX1 U2144 ( .A(n2323), .Y(n2263) );
  OR2X2 U2145 ( .A(n1793), .B(n1794), .Y(n2371) );
  INVX1 U2146 ( .A(n2371), .Y(n2264) );
  OR2X2 U2147 ( .A(n1791), .B(n1792), .Y(n2374) );
  INVX1 U2148 ( .A(n2374), .Y(n2265) );
  OR2X2 U2149 ( .A(SH[20]), .B(SH[24]), .Y(n2375) );
  INVX1 U2150 ( .A(n2375), .Y(n2266) );
  OR2X1 U2151 ( .A(n506), .B(n2418), .Y(n198) );
  INVX1 U2152 ( .A(n198), .Y(n2267) );
  OR2X1 U2153 ( .A(n507), .B(n2418), .Y(n199) );
  INVX1 U2154 ( .A(n199), .Y(n2268) );
  OR2X1 U2155 ( .A(n508), .B(n2418), .Y(n200) );
  INVX1 U2156 ( .A(n200), .Y(n2269) );
  OR2X1 U2157 ( .A(n509), .B(n2418), .Y(n201) );
  INVX1 U2158 ( .A(n201), .Y(n2270) );
  OR2X1 U2159 ( .A(n510), .B(n2418), .Y(n202) );
  INVX1 U2160 ( .A(n202), .Y(n2271) );
  OR2X1 U2161 ( .A(n515), .B(n2418), .Y(n207) );
  INVX1 U2162 ( .A(n207), .Y(n2272) );
  OR2X1 U2163 ( .A(n516), .B(n2418), .Y(n208) );
  INVX1 U2164 ( .A(n208), .Y(n2273) );
  OR2X1 U2165 ( .A(n517), .B(n2417), .Y(n209) );
  INVX1 U2166 ( .A(n209), .Y(n2274) );
  OR2X1 U2167 ( .A(n519), .B(n2417), .Y(n211) );
  INVX1 U2168 ( .A(n211), .Y(n2275) );
  OR2X1 U2169 ( .A(n520), .B(n2417), .Y(n212) );
  INVX1 U2170 ( .A(n212), .Y(n2276) );
  OR2X1 U2171 ( .A(n521), .B(n2417), .Y(n213) );
  INVX1 U2172 ( .A(n213), .Y(n2277) );
  OR2X1 U2173 ( .A(n522), .B(n2417), .Y(n214) );
  INVX1 U2174 ( .A(n214), .Y(n2278) );
  OR2X1 U2175 ( .A(n523), .B(n2417), .Y(n215) );
  INVX1 U2176 ( .A(n215), .Y(n2279) );
  INVX1 U2177 ( .A(n216), .Y(n2280) );
  OR2X1 U2178 ( .A(n525), .B(n2417), .Y(n217) );
  INVX1 U2179 ( .A(n217), .Y(n2281) );
  OR2X2 U2180 ( .A(n530), .B(n2417), .Y(n222) );
  INVX1 U2181 ( .A(n222), .Y(n2282) );
  OR2X2 U2182 ( .A(n531), .B(n2417), .Y(n223) );
  INVX1 U2183 ( .A(n223), .Y(n2283) );
  OR2X1 U2184 ( .A(n533), .B(n2417), .Y(n225) );
  INVX1 U2185 ( .A(n225), .Y(n2284) );
  OR2X1 U2186 ( .A(n535), .B(n2417), .Y(n227) );
  INVX1 U2187 ( .A(n227), .Y(n2285) );
  OR2X1 U2188 ( .A(n551), .B(n2416), .Y(n243) );
  INVX1 U2189 ( .A(n243), .Y(n2286) );
  OR2X2 U2190 ( .A(n553), .B(n2416), .Y(n245) );
  INVX1 U2191 ( .A(n245), .Y(n2287) );
  OR2X1 U2192 ( .A(n556), .B(n2416), .Y(n248) );
  INVX1 U2193 ( .A(n248), .Y(n2288) );
  OR2X1 U2194 ( .A(n564), .B(n2415), .Y(n256) );
  INVX1 U2195 ( .A(n256), .Y(n2289) );
  OR2X1 U2196 ( .A(n565), .B(n2415), .Y(n257) );
  INVX1 U2197 ( .A(n257), .Y(n2290) );
  OR2X2 U2198 ( .A(SH[28]), .B(SH[30]), .Y(n2324) );
  INVX1 U2199 ( .A(n2324), .Y(n2291) );
  INVX1 U2200 ( .A(n2376), .Y(n2292) );
  INVX1 U2201 ( .A(n2226), .Y(n2293) );
  INVX1 U2202 ( .A(n1782), .Y(n2294) );
  OR2X2 U2203 ( .A(n2398), .B(n711), .Y(n531) );
  OR2X1 U2204 ( .A(n513), .B(n2418), .Y(n205) );
  INVX1 U2205 ( .A(n205), .Y(n2295) );
  OR2X2 U2206 ( .A(n2399), .B(n693), .Y(n513) );
  OR2X2 U2207 ( .A(n2397), .B(n458), .Y(n545) );
  INVX1 U2208 ( .A(n2245), .Y(n2296) );
  INVX1 U2209 ( .A(n2296), .Y(n2297) );
  INVX1 U2210 ( .A(n2248), .Y(n2298) );
  INVX1 U2211 ( .A(n2298), .Y(n2299) );
  INVX1 U2212 ( .A(n2253), .Y(n2300) );
  INVX1 U2213 ( .A(n2300), .Y(n2301) );
  AND2X2 U2214 ( .A(n307), .B(n2333), .Y(B[113]) );
  OR2X2 U2215 ( .A(n2399), .B(n687), .Y(n507) );
  OR2X2 U2216 ( .A(n538), .B(n2416), .Y(n230) );
  INVX1 U2217 ( .A(n230), .Y(n2302) );
  OR2X2 U2218 ( .A(n2397), .B(n465), .Y(n538) );
  OR2X2 U2219 ( .A(n546), .B(n2416), .Y(n238) );
  INVX1 U2220 ( .A(n238), .Y(n2303) );
  OR2X2 U2221 ( .A(n2397), .B(n457), .Y(n546) );
  OR2X2 U2222 ( .A(n547), .B(n2416), .Y(n239) );
  INVX1 U2223 ( .A(n239), .Y(n2304) );
  OR2X2 U2224 ( .A(n2397), .B(n456), .Y(n547) );
  OR2X2 U2225 ( .A(n548), .B(n2416), .Y(n240) );
  INVX1 U2226 ( .A(n240), .Y(n2305) );
  OR2X2 U2227 ( .A(n2397), .B(n455), .Y(n548) );
  OR2X2 U2228 ( .A(n549), .B(n2416), .Y(n241) );
  INVX1 U2229 ( .A(n241), .Y(n2306) );
  OR2X2 U2230 ( .A(n2397), .B(n454), .Y(n549) );
  OR2X2 U2231 ( .A(n534), .B(n2417), .Y(n226) );
  INVX1 U2232 ( .A(n226), .Y(n2307) );
  AND2X2 U2233 ( .A(n283), .B(n2379), .Y(B[89]) );
  AND2X2 U2234 ( .A(n309), .B(n2384), .Y(B[115]) );
  AND2X2 U2235 ( .A(n359), .B(n2316), .Y(B[165]) );
  AND2X2 U2236 ( .A(n371), .B(n2333), .Y(B[177]) );
  AND2X2 U2237 ( .A(n339), .B(n2383), .Y(B[145]) );
  INVX1 U2238 ( .A(n2322), .Y(n2308) );
  INVX1 U2239 ( .A(n683), .Y(n2309) );
  INVX1 U2240 ( .A(n684), .Y(n2310) );
  OR2X2 U2241 ( .A(n2462), .B(n1060), .Y(n880) );
  INVX1 U2242 ( .A(n685), .Y(n2311) );
  OR2X2 U2243 ( .A(n888), .B(n2439), .Y(n692) );
  INVX1 U2244 ( .A(n692), .Y(n2312) );
  OR2X2 U2245 ( .A(n2461), .B(n867), .Y(n888) );
  INVX1 U2246 ( .A(n693), .Y(n2313) );
  INVX1 U2247 ( .A(n709), .Y(n2314) );
  AND2X2 U2248 ( .A(n311), .B(n2318), .Y(B[117]) );
  AND2X2 U2249 ( .A(n351), .B(n2316), .Y(B[157]) );
  AND2X2 U2250 ( .A(n292), .B(n2315), .Y(B[98]) );
  AND2X2 U2251 ( .A(n294), .B(n2384), .Y(B[100]) );
  AND2X2 U2252 ( .A(n296), .B(n2381), .Y(B[102]) );
  AND2X2 U2253 ( .A(n298), .B(n2315), .Y(B[104]) );
  AND2X2 U2254 ( .A(n300), .B(n2315), .Y(B[106]) );
  AND2X2 U2255 ( .A(n302), .B(n2223), .Y(B[108]) );
  AND2X2 U2256 ( .A(n304), .B(n2315), .Y(B[110]) );
  AND2X2 U2257 ( .A(n306), .B(n2318), .Y(B[112]) );
  AND2X2 U2258 ( .A(n316), .B(n2318), .Y(B[122]) );
  AND2X2 U2259 ( .A(n318), .B(n2381), .Y(B[124]) );
  AND2X2 U2260 ( .A(n322), .B(n2384), .Y(B[128]) );
  AND2X2 U2261 ( .A(n342), .B(n2381), .Y(B[148]) );
  AND2X2 U2262 ( .A(n360), .B(n2382), .Y(B[166]) );
  AND2X2 U2263 ( .A(n362), .B(n2384), .Y(B[168]) );
  AND2X2 U2264 ( .A(n277), .B(n2381), .Y(B[83]) );
  AND2X2 U2265 ( .A(n279), .B(n2315), .Y(B[85]) );
  AND2X2 U2266 ( .A(n281), .B(n2381), .Y(B[87]) );
  AND2X2 U2267 ( .A(n287), .B(n2381), .Y(B[93]) );
  AND2X2 U2268 ( .A(n291), .B(n2383), .Y(B[97]) );
  AND2X2 U2269 ( .A(n295), .B(n2384), .Y(B[101]) );
  AND2X2 U2270 ( .A(n297), .B(n2380), .Y(B[103]) );
  AND2X2 U2271 ( .A(n301), .B(n2331), .Y(B[107]) );
  AND2X2 U2272 ( .A(n303), .B(n2384), .Y(B[109]) );
  AND2X2 U2273 ( .A(n337), .B(n2316), .Y(B[143]) );
  AND2X2 U2274 ( .A(n341), .B(n2384), .Y(B[147]) );
  AND2X2 U2275 ( .A(n345), .B(n2384), .Y(B[151]) );
  AND2X2 U2276 ( .A(n357), .B(n2315), .Y(B[163]) );
  AND2X2 U2277 ( .A(n365), .B(n2223), .Y(B[171]) );
  AND2X2 U2278 ( .A(n369), .B(n2315), .Y(B[175]) );
  AND2X2 U2279 ( .A(n290), .B(n2318), .Y(B[96]) );
  AND2X2 U2280 ( .A(n314), .B(n2315), .Y(B[120]) );
  AND2X2 U2281 ( .A(n338), .B(n2333), .Y(B[144]) );
  AND2X2 U2282 ( .A(n346), .B(n2315), .Y(B[152]) );
  AND2X2 U2283 ( .A(n348), .B(n2318), .Y(B[154]) );
  AND2X2 U2284 ( .A(n352), .B(n2384), .Y(B[158]) );
  AND2X2 U2285 ( .A(n354), .B(n2382), .Y(B[160]) );
  AND2X2 U2286 ( .A(n356), .B(n2384), .Y(B[162]) );
  AND2X2 U2287 ( .A(n358), .B(n2384), .Y(B[164]) );
  AND2X2 U2288 ( .A(n364), .B(n2381), .Y(B[170]) );
  AND2X2 U2289 ( .A(n366), .B(n2384), .Y(B[172]) );
  AND2X2 U2290 ( .A(n368), .B(n2381), .Y(B[174]) );
  AND2X2 U2291 ( .A(n370), .B(n2384), .Y(B[176]) );
  OR2X2 U2292 ( .A(SH[27]), .B(SH[25]), .Y(n1793) );
  OR2X2 U2293 ( .A(n884), .B(n2439), .Y(n688) );
  OR2X2 U2294 ( .A(n2500), .B(n1422), .Y(n1242) );
  INVX2 U2295 ( .A(SH[2]), .Y(n2502) );
  OR2X2 U2296 ( .A(n2398), .B(n699), .Y(n519) );
  INVX4 U2297 ( .A(n2502), .Y(n2496) );
  INVX4 U2298 ( .A(n2317), .Y(n2318) );
  INVX2 U2299 ( .A(n2446), .Y(n2466) );
  INVX8 U2300 ( .A(n2483), .Y(n2468) );
  INVX1 U2301 ( .A(n1782), .Y(n2317) );
  INVX4 U2302 ( .A(n2482), .Y(n2474) );
  OR2X2 U2303 ( .A(n2500), .B(n1240), .Y(n1243) );
  INVX2 U2304 ( .A(SH[1]), .Y(n2507) );
  INVX2 U2305 ( .A(n2525), .Y(n2519) );
  OR2X2 U2306 ( .A(n2399), .B(n688), .Y(n508) );
  INVX4 U2307 ( .A(n2226), .Y(n2386) );
  OR2X2 U2308 ( .A(n1243), .B(n2208), .Y(n879) );
  INVX4 U2309 ( .A(n2506), .Y(n2525) );
  OR2X2 U2310 ( .A(n2462), .B(n874), .Y(n881) );
  INVX2 U2311 ( .A(n2525), .Y(n2515) );
  INVX1 U2312 ( .A(n2525), .Y(n2321) );
  INVX2 U2313 ( .A(n2400), .Y(n2397) );
  OR2X2 U2314 ( .A(n2399), .B(n689), .Y(n509) );
  OR2X2 U2315 ( .A(n1801), .B(n1802), .Y(n1791) );
  AND2X2 U2316 ( .A(n289), .B(n2379), .Y(B[95]) );
  AND2X2 U2317 ( .A(n2263), .B(n2291), .Y(n2377) );
  INVX2 U2318 ( .A(n2482), .Y(n2480) );
  INVX4 U2319 ( .A(n2501), .Y(n2495) );
  BUFX4 U2320 ( .A(n2477), .Y(n2325) );
  INVX4 U2321 ( .A(n2481), .Y(n2477) );
  INVX2 U2322 ( .A(n2477), .Y(n2483) );
  AND2X2 U2323 ( .A(n285), .B(n2381), .Y(B[91]) );
  OR2X1 U2324 ( .A(n502), .B(n2418), .Y(n194) );
  INVX1 U2325 ( .A(n2226), .Y(n2385) );
  AND2X2 U2326 ( .A(n350), .B(n2384), .Y(B[156]) );
  INVX1 U2327 ( .A(n2478), .Y(n2328) );
  OR2X2 U2328 ( .A(n2396), .B(n435), .Y(n568) );
  AND2X2 U2329 ( .A(n2373), .B(n2265), .Y(n2327) );
  OR2X2 U2330 ( .A(SH[14]), .B(SH[12]), .Y(n1802) );
  AND2X2 U2331 ( .A(n344), .B(n2223), .Y(B[150]) );
  INVX1 U2332 ( .A(n2485), .Y(n2326) );
  INVX2 U2333 ( .A(SH[2]), .Y(n2485) );
  MUX2X1 U2334 ( .B(n1264), .A(n1272), .S(n2328), .Y(n1088) );
  MUX2X1 U2335 ( .B(n1700), .A(n1702), .S(n2525), .Y(n1522) );
  MUX2X1 U2336 ( .B(n1148), .A(n1164), .S(n2334), .Y(n984) );
  AND2X2 U2337 ( .A(n340), .B(n2384), .Y(B[146]) );
  AND2X2 U2338 ( .A(n293), .B(n2318), .Y(B[99]) );
  AND2X2 U2339 ( .A(n305), .B(n2316), .Y(B[111]) );
  AND2X2 U2340 ( .A(n2258), .B(n2384), .Y(B[58]) );
  AND2X2 U2341 ( .A(n2260), .B(n2384), .Y(B[60]) );
  AND2X2 U2342 ( .A(n2268), .B(n2384), .Y(B[5]) );
  INVX1 U2343 ( .A(n1300), .Y(n2329) );
  INVX1 U2344 ( .A(n2329), .Y(n2330) );
  INVX8 U2345 ( .A(n2386), .Y(n2384) );
  INVX2 U2346 ( .A(n2485), .Y(n2500) );
  INVX4 U2347 ( .A(n2443), .Y(n2429) );
  INVX4 U2348 ( .A(n2482), .Y(n2471) );
  INVX4 U2349 ( .A(n2482), .Y(n2475) );
  INVX4 U2350 ( .A(n2482), .Y(n2476) );
  INVX4 U2351 ( .A(n2482), .Y(n2470) );
  AND2X2 U2352 ( .A(n336), .B(n2316), .Y(B[142]) );
  INVX4 U2353 ( .A(n2465), .Y(n2451) );
  INVX1 U2354 ( .A(n460), .Y(n2332) );
  AND2X2 U2355 ( .A(n310), .B(n2381), .Y(B[116]) );
  OR2X2 U2356 ( .A(n2461), .B(n866), .Y(n889) );
  AND2X2 U2357 ( .A(n320), .B(n2333), .Y(B[126]) );
  MUX2X1 U2358 ( .B(n1106), .A(n1122), .S(n2466), .Y(n942) );
  AND2X2 U2359 ( .A(n334), .B(n2381), .Y(B[140]) );
  MUX2X1 U2360 ( .B(n1140), .A(n1156), .S(n2334), .Y(n976) );
  INVX4 U2361 ( .A(n2464), .Y(n2454) );
  INVX2 U2362 ( .A(n2461), .Y(n2334) );
  INVX4 U2363 ( .A(n2502), .Y(n2493) );
  AND2X2 U2364 ( .A(n312), .B(n2333), .Y(B[118]) );
  OR2X2 U2365 ( .A(n2399), .B(n691), .Y(n511) );
  AND2X2 U2366 ( .A(n2235), .B(n2381), .Y(B[10]) );
  INVX4 U2367 ( .A(n2443), .Y(n2428) );
  AND2X2 U2368 ( .A(n2270), .B(n2379), .Y(B[7]) );
  OR2X2 U2369 ( .A(n2396), .B(n437), .Y(n566) );
  MUX2X1 U2370 ( .B(n1100), .A(n1116), .S(n2466), .Y(n936) );
  MUX2X1 U2371 ( .B(n1620), .A(n1622), .S(n2525), .Y(n1442) );
  INVX2 U2372 ( .A(n2523), .Y(n2521) );
  INVX2 U2373 ( .A(n2523), .Y(n2520) );
  MUX2X1 U2374 ( .B(n1644), .A(n1646), .S(n2525), .Y(n1466) );
  AND2X2 U2375 ( .A(n330), .B(n2384), .Y(B[136]) );
  AND2X2 U2376 ( .A(n328), .B(n2384), .Y(B[134]) );
  AND2X2 U2377 ( .A(n308), .B(n2380), .Y(B[114]) );
  AND2X2 U2378 ( .A(n326), .B(n2221), .Y(B[132]) );
  INVX8 U2379 ( .A(n2444), .Y(n2426) );
  OR2X2 U2380 ( .A(n878), .B(n2439), .Y(n2335) );
  OR2X2 U2381 ( .A(n2462), .B(n2322), .Y(n878) );
  INVX4 U2382 ( .A(n2440), .Y(n2439) );
  MUX2X1 U2383 ( .B(n1654), .A(n1656), .S(n2525), .Y(n1476) );
  AND2X2 U2384 ( .A(n282), .B(n2316), .Y(B[88]) );
  AND2X2 U2385 ( .A(n278), .B(n2221), .Y(B[84]) );
  MUX2X1 U2386 ( .B(n934), .A(n966), .S(n2444), .Y(n770) );
  INVX2 U2387 ( .A(n2442), .Y(n2433) );
  MUX2X1 U2388 ( .B(n1438), .A(n1442), .S(n2504), .Y(n1262) );
  INVX2 U2389 ( .A(n2484), .Y(n2504) );
  AND2X2 U2390 ( .A(n332), .B(n2382), .Y(B[138]) );
  MUX2X1 U2391 ( .B(n1612), .A(n1614), .S(n2525), .Y(n1434) );
  INVX2 U2392 ( .A(n2502), .Y(n2494) );
  AND2X2 U2393 ( .A(n324), .B(n2379), .Y(B[130]) );
  INVX2 U2394 ( .A(n2482), .Y(n2473) );
  INVX2 U2395 ( .A(n2482), .Y(n2472) );
  INVX2 U2396 ( .A(n2481), .Y(n2478) );
  OR2X2 U2397 ( .A(n1249), .B(n2471), .Y(n1065) );
  OR2X2 U2398 ( .A(n1246), .B(n2475), .Y(n1062) );
  OR2X2 U2399 ( .A(n1248), .B(n2480), .Y(n1064) );
  OR2X2 U2400 ( .A(n1247), .B(n2471), .Y(n1063) );
  INVX2 U2401 ( .A(n2294), .Y(n2379) );
  MUX2X1 U2402 ( .B(n1436), .A(n1440), .S(n2504), .Y(n1260) );
  AND2X2 U2403 ( .A(n2282), .B(n2318), .Y(B[28]) );
  AND2X2 U2404 ( .A(n2240), .B(n2318), .Y(B[26]) );
  AND2X2 U2405 ( .A(n2238), .B(n2318), .Y(B[24]) );
  AND2X2 U2406 ( .A(n2281), .B(n2318), .Y(B[23]) );
  AND2X2 U2407 ( .A(n2279), .B(n2381), .Y(B[21]) );
  AND2X2 U2408 ( .A(n2277), .B(n2380), .Y(B[19]) );
  AND2X2 U2409 ( .A(n2267), .B(n2379), .Y(B[4]) );
  AND2X2 U2410 ( .A(n2236), .B(n2333), .Y(B[12]) );
  AND2X2 U2411 ( .A(n361), .B(n2223), .Y(B[167]) );
  AND2X2 U2412 ( .A(n363), .B(n2223), .Y(B[169]) );
  AND2X2 U2413 ( .A(n367), .B(n2384), .Y(B[173]) );
  AND2X2 U2414 ( .A(n2288), .B(n2381), .Y(B[54]) );
  AND2X2 U2415 ( .A(n372), .B(n2315), .Y(B[178]) );
  AND2X2 U2416 ( .A(n2304), .B(n2333), .Y(B[45]) );
  AND2X2 U2417 ( .A(n2302), .B(n2333), .Y(B[36]) );
  AND2X2 U2418 ( .A(n2246), .B(n2381), .Y(B[38]) );
  AND2X2 U2419 ( .A(n2287), .B(n2379), .Y(B[51]) );
  AND2X2 U2420 ( .A(n2254), .B(n2333), .Y(B[53]) );
  AND2X2 U2421 ( .A(n2306), .B(n2316), .Y(B[47]) );
  AND2X2 U2422 ( .A(n2286), .B(n2384), .Y(B[49]) );
  AND2X2 U2423 ( .A(n2250), .B(n2333), .Y(B[42]) );
  AND2X2 U2424 ( .A(n2256), .B(n2384), .Y(B[56]) );
  INVX2 U2425 ( .A(n2441), .Y(n2434) );
  AND2X2 U2426 ( .A(n2242), .B(n2318), .Y(B[30]) );
  AND2X2 U2427 ( .A(n280), .B(n2221), .Y(B[86]) );
  INVX2 U2428 ( .A(n2502), .Y(n2498) );
  AND2X2 U2429 ( .A(n274), .B(n2316), .Y(B[80]) );
  INVX2 U2430 ( .A(n2485), .Y(n2497) );
  AND2X2 U2431 ( .A(n2233), .B(n2318), .Y(B[3]) );
  AND2X2 U2432 ( .A(n2231), .B(n2225), .Y(B[1]) );
  AND2X2 U2433 ( .A(n2232), .B(n2225), .Y(B[2]) );
  AND2X2 U2434 ( .A(n276), .B(n2381), .Y(B[82]) );
  AND2X2 U2435 ( .A(n2274), .B(n2318), .Y(B[15]) );
  INVX2 U2436 ( .A(SH[4]), .Y(n2447) );
  AND2X2 U2437 ( .A(n2383), .B(n2234), .Y(B[9]) );
  AND2X2 U2438 ( .A(n2271), .B(n2318), .Y(B[8]) );
  INVX2 U2439 ( .A(n2442), .Y(n2336) );
  INVX2 U2440 ( .A(n2442), .Y(n2337) );
  INVX4 U2441 ( .A(n2464), .Y(n2456) );
  INVX4 U2442 ( .A(n2464), .Y(n2455) );
  AND2X2 U2443 ( .A(n270), .B(n2333), .Y(B[76]) );
  AND2X2 U2444 ( .A(n288), .B(n2315), .Y(B[94]) );
  AND2X2 U2445 ( .A(n286), .B(n2382), .Y(B[92]) );
  AND2X2 U2446 ( .A(n264), .B(n2381), .Y(B[70]) );
  AND2X2 U2447 ( .A(n262), .B(n2331), .Y(B[68]) );
  INVX2 U2448 ( .A(SH[3]), .Y(n2481) );
  INVX2 U2449 ( .A(SH[3]), .Y(n2482) );
  MUX2X1 U2450 ( .B(n1104), .A(n1120), .S(n2466), .Y(n940) );
  INVX1 U2451 ( .A(n2447), .Y(n2457) );
  AND2X2 U2452 ( .A(n272), .B(n2379), .Y(B[78]) );
  AND2X2 U2453 ( .A(n284), .B(n2221), .Y(B[90]) );
  OR2X2 U2454 ( .A(n2394), .B(n407), .Y(n596) );
  OR2X2 U2455 ( .A(n411), .B(n2395), .Y(n592) );
  OR2X2 U2456 ( .A(n2398), .B(n708), .Y(n528) );
  OR2X1 U2457 ( .A(n887), .B(n2439), .Y(n691) );
  AND2X2 U2458 ( .A(n333), .B(n2384), .Y(B[139]) );
  AND2X2 U2459 ( .A(n335), .B(n2315), .Y(B[141]) );
  AND2X2 U2460 ( .A(n331), .B(n2223), .Y(B[137]) );
  AND2X2 U2461 ( .A(n329), .B(n2384), .Y(B[135]) );
  AND2X2 U2462 ( .A(n327), .B(n2333), .Y(B[133]) );
  AND2X2 U2463 ( .A(n321), .B(n2316), .Y(B[127]) );
  AND2X2 U2464 ( .A(n325), .B(n2315), .Y(B[131]) );
  AND2X2 U2465 ( .A(n317), .B(n2316), .Y(B[123]) );
  AND2X2 U2466 ( .A(n323), .B(n2381), .Y(B[129]) );
  AND2X2 U2467 ( .A(n2289), .B(n2384), .Y(B[62]) );
  AND2X2 U2468 ( .A(n315), .B(n2315), .Y(B[121]) );
  AND2X2 U2469 ( .A(n319), .B(n2315), .Y(B[125]) );
  AND2X2 U2470 ( .A(n313), .B(n2384), .Y(B[119]) );
  AND2X2 U2471 ( .A(n2295), .B(n2384), .Y(B[11]) );
  AND2X2 U2472 ( .A(n2272), .B(n2223), .Y(B[13]) );
  OR2X2 U2473 ( .A(n2399), .B(n690), .Y(n510) );
  AND2X2 U2474 ( .A(n2299), .B(n2221), .Y(B[40]) );
  OR2X2 U2475 ( .A(n2398), .B(n469), .Y(n534) );
  AND2X2 U2476 ( .A(n373), .B(n2384), .Y(B[179]) );
  AND2X2 U2477 ( .A(n2305), .B(n2315), .Y(B[46]) );
  AND2X2 U2478 ( .A(n2257), .B(n2333), .Y(B[57]) );
  AND2X2 U2479 ( .A(n2303), .B(n2315), .Y(B[44]) );
  AND2X2 U2480 ( .A(n2255), .B(n2331), .Y(B[55]) );
  AND2X2 U2481 ( .A(n2249), .B(n2381), .Y(B[41]) );
  AND2X2 U2482 ( .A(n266), .B(n2333), .Y(B[72]) );
  AND2X2 U2483 ( .A(n2301), .B(n2384), .Y(B[50]) );
  AND2X2 U2484 ( .A(n2297), .B(n2382), .Y(B[37]) );
  AND2X2 U2485 ( .A(n2247), .B(n2381), .Y(B[39]) );
  AND2X2 U2486 ( .A(n2252), .B(n2331), .Y(B[48]) );
  AND2X2 U2487 ( .A(n2228), .B(n2318), .Y(B[52]) );
  AND2X2 U2488 ( .A(n260), .B(n2331), .Y(B[66]) );
  AND2X2 U2489 ( .A(n273), .B(n2315), .Y(B[79]) );
  AND2X2 U2490 ( .A(n269), .B(n2333), .Y(B[75]) );
  AND2X2 U2491 ( .A(n271), .B(n2316), .Y(B[77]) );
  AND2X2 U2492 ( .A(n267), .B(n2331), .Y(B[73]) );
  AND2X2 U2493 ( .A(n2261), .B(n2333), .Y(B[61]) );
  AND2X2 U2494 ( .A(n265), .B(n2380), .Y(B[71]) );
  AND2X2 U2495 ( .A(n2290), .B(n2333), .Y(B[63]) );
  AND2X2 U2496 ( .A(n275), .B(n2333), .Y(B[81]) );
  AND2X2 U2497 ( .A(n263), .B(n2380), .Y(B[69]) );
  AND2X2 U2498 ( .A(n261), .B(n2380), .Y(B[67]) );
  AND2X2 U2499 ( .A(n2259), .B(n2381), .Y(B[59]) );
  AND2X2 U2500 ( .A(n259), .B(n2331), .Y(B[65]) );
  AND2X2 U2501 ( .A(n258), .B(n2315), .Y(B[64]) );
  OR2X2 U2502 ( .A(n899), .B(n2438), .Y(n703) );
  INVX1 U2503 ( .A(n703), .Y(n2338) );
  OR2X2 U2504 ( .A(n885), .B(n2439), .Y(n689) );
  INVX1 U2505 ( .A(n689), .Y(n2339) );
  OR2X2 U2506 ( .A(n2462), .B(n1065), .Y(n885) );
  OR2X2 U2507 ( .A(n904), .B(n2438), .Y(n708) );
  INVX1 U2508 ( .A(n708), .Y(n2340) );
  OR2X2 U2509 ( .A(n895), .B(n2439), .Y(n699) );
  INVX1 U2510 ( .A(n699), .Y(n2341) );
  OR2X2 U2511 ( .A(n909), .B(n2438), .Y(n713) );
  INVX1 U2512 ( .A(n713), .Y(n2342) );
  OR2X1 U2513 ( .A(n883), .B(n2439), .Y(n687) );
  INVX1 U2514 ( .A(n687), .Y(n2343) );
  OR2X2 U2515 ( .A(n2462), .B(n1063), .Y(n883) );
  OR2X2 U2516 ( .A(n903), .B(n2438), .Y(n707) );
  INVX1 U2517 ( .A(n707), .Y(n2344) );
  OR2X2 U2518 ( .A(n893), .B(n2439), .Y(n697) );
  INVX1 U2519 ( .A(n697), .Y(n2345) );
  OR2X2 U2520 ( .A(n2461), .B(n862), .Y(n893) );
  OR2X2 U2521 ( .A(n2475), .B(n1245), .Y(n1061) );
  INVX1 U2522 ( .A(n1061), .Y(n2346) );
  INVX1 U2523 ( .A(n1061), .Y(n2347) );
  OR2X2 U2524 ( .A(n901), .B(n2438), .Y(n705) );
  INVX1 U2525 ( .A(n705), .Y(n2348) );
  OR2X2 U2526 ( .A(n894), .B(n2439), .Y(n698) );
  INVX1 U2527 ( .A(n698), .Y(n2349) );
  OR2X2 U2528 ( .A(n2471), .B(n1244), .Y(n1060) );
  INVX1 U2529 ( .A(n1060), .Y(n2350) );
  OR2X2 U2530 ( .A(n907), .B(n2438), .Y(n711) );
  INVX1 U2531 ( .A(n711), .Y(n2351) );
  INVX1 U2532 ( .A(n691), .Y(n2352) );
  OR2X2 U2533 ( .A(n2461), .B(n868), .Y(n887) );
  OR2X2 U2534 ( .A(n2480), .B(n1243), .Y(n1059) );
  OR2X2 U2535 ( .A(n896), .B(n2438), .Y(n700) );
  INVX1 U2536 ( .A(n700), .Y(n2353) );
  OR2X2 U2537 ( .A(n892), .B(n2439), .Y(n696) );
  INVX1 U2538 ( .A(n696), .Y(n2354) );
  OR2X2 U2539 ( .A(n2461), .B(n863), .Y(n892) );
  OR2X2 U2540 ( .A(n908), .B(n2438), .Y(n712) );
  INVX1 U2541 ( .A(n712), .Y(n2355) );
  OR2X2 U2542 ( .A(n891), .B(n2439), .Y(n695) );
  INVX1 U2543 ( .A(n695), .Y(n2356) );
  OR2X2 U2544 ( .A(n2461), .B(n864), .Y(n891) );
  OR2X2 U2545 ( .A(n898), .B(n2438), .Y(n702) );
  INVX1 U2546 ( .A(n702), .Y(n2357) );
  INVX1 U2547 ( .A(n1065), .Y(n2358) );
  INVX1 U2548 ( .A(n688), .Y(n2359) );
  OR2X2 U2549 ( .A(n2462), .B(n1064), .Y(n884) );
  OR2X2 U2550 ( .A(n906), .B(n2438), .Y(n710) );
  INVX1 U2551 ( .A(n710), .Y(n2360) );
  INVX1 U2552 ( .A(n1064), .Y(n2361) );
  OR2X2 U2553 ( .A(n890), .B(n2439), .Y(n694) );
  INVX1 U2554 ( .A(n694), .Y(n2362) );
  OR2X2 U2555 ( .A(n2461), .B(n865), .Y(n890) );
  INVX1 U2556 ( .A(n194), .Y(n2363) );
  OR2X2 U2557 ( .A(n2399), .B(n2335), .Y(n502) );
  OR2X2 U2558 ( .A(n2522), .B(n1602), .Y(n1422) );
  OR2X2 U2559 ( .A(n902), .B(n2438), .Y(n706) );
  INVX1 U2560 ( .A(n706), .Y(n2365) );
  OR2X1 U2561 ( .A(n882), .B(n2439), .Y(n686) );
  INVX1 U2562 ( .A(n686), .Y(n2366) );
  OR2X2 U2563 ( .A(n2462), .B(n1062), .Y(n882) );
  AND2X2 U2564 ( .A(n2264), .B(n2372), .Y(n1784) );
  OR2X2 U2565 ( .A(n1603), .B(n2522), .Y(n1423) );
  INVX1 U2566 ( .A(n1423), .Y(n2367) );
  INVX1 U2567 ( .A(n1423), .Y(n2368) );
  OR2X2 U2568 ( .A(n900), .B(n2438), .Y(n704) );
  INVX1 U2569 ( .A(n704), .Y(n2369) );
  OR2X1 U2570 ( .A(n886), .B(n2439), .Y(n690) );
  INVX1 U2571 ( .A(n690), .Y(n2370) );
  OR2X2 U2572 ( .A(n2462), .B(n869), .Y(n886) );
  INVX2 U2573 ( .A(n2441), .Y(n2435) );
  INVX2 U2574 ( .A(n2419), .Y(n2416) );
  INVX2 U2575 ( .A(n2503), .Y(n2491) );
  INVX1 U2576 ( .A(n2421), .Y(n2412) );
  INVX2 U2577 ( .A(n2503), .Y(n2490) );
  INVX2 U2578 ( .A(n2443), .Y(n2430) );
  INVX2 U2579 ( .A(n2524), .Y(n2512) );
  INVX1 U2580 ( .A(n2222), .Y(n2382) );
  INVX2 U2581 ( .A(n2402), .Y(n2393) );
  INVX2 U2582 ( .A(n2400), .Y(n2398) );
  INVX2 U2583 ( .A(n2401), .Y(n2396) );
  INVX2 U2584 ( .A(n2419), .Y(n2417) );
  INVX2 U2585 ( .A(n2420), .Y(n2415) );
  INVX2 U2586 ( .A(n2463), .Y(n2460) );
  INVX2 U2587 ( .A(n2465), .Y(n2452) );
  INVX2 U2588 ( .A(n2465), .Y(n2453) );
  INVX2 U2589 ( .A(n2504), .Y(n2487) );
  INVX2 U2590 ( .A(n2504), .Y(n2488) );
  INVX2 U2591 ( .A(n2483), .Y(n2467) );
  INVX2 U2592 ( .A(n2466), .Y(n2449) );
  INVX2 U2593 ( .A(n2466), .Y(n2450) );
  INVX2 U2594 ( .A(n2444), .Y(n2427) );
  INVX2 U2595 ( .A(n2524), .Y(n2513) );
  INVX2 U2596 ( .A(n2525), .Y(n2509) );
  INVX2 U2597 ( .A(n2525), .Y(n2510) );
  INVX2 U2598 ( .A(n2402), .Y(n2390) );
  OR2X2 U2599 ( .A(n1803), .B(SH[29]), .Y(n1792) );
  INVX1 U2600 ( .A(SH[5]), .Y(n2425) );
  INVX1 U2601 ( .A(SH[7]), .Y(n2388) );
  INVX1 U2602 ( .A(SH[6]), .Y(n2405) );
  INVX1 U2603 ( .A(n2222), .Y(n2383) );
  INVX1 U2604 ( .A(n803), .Y(n380) );
  INVX1 U2605 ( .A(n799), .Y(n384) );
  INVX1 U2606 ( .A(n801), .Y(n382) );
  INVX1 U2607 ( .A(n807), .Y(n376) );
  INVX1 U2608 ( .A(n805), .Y(n378) );
  INVX1 U2609 ( .A(n809), .Y(n374) );
  INVX1 U2610 ( .A(n802), .Y(n381) );
  INVX1 U2611 ( .A(n798), .Y(n385) );
  INVX1 U2612 ( .A(n800), .Y(n383) );
  INVX1 U2613 ( .A(n806), .Y(n377) );
  INVX1 U2614 ( .A(n804), .Y(n379) );
  INVX1 U2615 ( .A(n808), .Y(n375) );
  INVX1 U2616 ( .A(n776), .Y(n407) );
  INVX1 U2617 ( .A(n774), .Y(n409) );
  INVX1 U2618 ( .A(n778), .Y(n405) );
  INVX1 U2619 ( .A(n772), .Y(n411) );
  INVX1 U2620 ( .A(n770), .Y(n413) );
  INVX1 U2621 ( .A(n764), .Y(n419) );
  INVX1 U2622 ( .A(n750), .Y(n433) );
  INVX1 U2623 ( .A(n748), .Y(n435) );
  INVX1 U2624 ( .A(n780), .Y(n403) );
  INVX1 U2625 ( .A(n768), .Y(n415) );
  INVX1 U2626 ( .A(n762), .Y(n421) );
  INVX1 U2627 ( .A(n754), .Y(n429) );
  INVX1 U2628 ( .A(n766), .Y(n417) );
  INVX1 U2629 ( .A(n760), .Y(n423) );
  INVX1 U2630 ( .A(n794), .Y(n389) );
  INVX1 U2631 ( .A(n752), .Y(n431) );
  INVX1 U2632 ( .A(n792), .Y(n391) );
  INVX1 U2633 ( .A(n777), .Y(n406) );
  INVX1 U2634 ( .A(n786), .Y(n397) );
  INVX1 U2635 ( .A(n756), .Y(n427) );
  INVX1 U2636 ( .A(n758), .Y(n425) );
  INVX1 U2637 ( .A(n782), .Y(n401) );
  INVX1 U2638 ( .A(n775), .Y(n408) );
  INVX1 U2639 ( .A(n788), .Y(n395) );
  INVX1 U2640 ( .A(n790), .Y(n393) );
  INVX1 U2641 ( .A(n784), .Y(n399) );
  INVX1 U2642 ( .A(n746), .Y(n437) );
  INVX1 U2643 ( .A(n779), .Y(n404) );
  INVX1 U2644 ( .A(n747), .Y(n436) );
  INVX1 U2645 ( .A(n793), .Y(n390) );
  INVX1 U2646 ( .A(n773), .Y(n410) );
  INVX1 U2647 ( .A(n761), .Y(n422) );
  INVX1 U2648 ( .A(n763), .Y(n420) );
  INVX1 U2649 ( .A(n749), .Y(n434) );
  INVX1 U2650 ( .A(n795), .Y(n388) );
  INVX1 U2651 ( .A(n781), .Y(n402) );
  INVX1 U2652 ( .A(n751), .Y(n432) );
  INVX1 U2653 ( .A(n771), .Y(n412) );
  INVX1 U2654 ( .A(n755), .Y(n428) );
  INVX1 U2655 ( .A(n765), .Y(n418) );
  INVX1 U2656 ( .A(n769), .Y(n414) );
  INVX1 U2657 ( .A(n787), .Y(n396) );
  INVX1 U2658 ( .A(n759), .Y(n424) );
  INVX1 U2659 ( .A(n767), .Y(n416) );
  INVX1 U2660 ( .A(n753), .Y(n430) );
  INVX1 U2661 ( .A(n757), .Y(n426) );
  INVX1 U2662 ( .A(n789), .Y(n394) );
  INVX1 U2663 ( .A(n783), .Y(n400) );
  INVX1 U2664 ( .A(n791), .Y(n392) );
  INVX1 U2665 ( .A(n785), .Y(n398) );
  INVX1 U2666 ( .A(n796), .Y(n387) );
  INVX1 U2667 ( .A(n797), .Y(n386) );
  INVX1 U2668 ( .A(n728), .Y(n455) );
  INVX1 U2669 ( .A(n729), .Y(n454) );
  INVX1 U2670 ( .A(n736), .Y(n447) );
  INVX1 U2671 ( .A(n730), .Y(n453) );
  INVX1 U2672 ( .A(n732), .Y(n451) );
  INVX1 U2673 ( .A(n738), .Y(n445) );
  INVX1 U2674 ( .A(n716), .Y(n467) );
  INVX1 U2675 ( .A(n726), .Y(n457) );
  INVX1 U2676 ( .A(n718), .Y(n465) );
  INVX1 U2677 ( .A(n734), .Y(n449) );
  INVX1 U2678 ( .A(n724), .Y(n459) );
  INVX1 U2679 ( .A(n737), .Y(n446) );
  INVX1 U2680 ( .A(n720), .Y(n463) );
  INVX1 U2681 ( .A(n744), .Y(n439) );
  INVX1 U2682 ( .A(n742), .Y(n441) );
  INVX1 U2683 ( .A(n731), .Y(n452) );
  INVX1 U2684 ( .A(n740), .Y(n443) );
  INVX1 U2685 ( .A(n717), .Y(n466) );
  INVX1 U2686 ( .A(n727), .Y(n456) );
  INVX1 U2687 ( .A(n739), .Y(n444) );
  INVX1 U2688 ( .A(n719), .Y(n464) );
  INVX1 U2689 ( .A(n733), .Y(n450) );
  INVX1 U2690 ( .A(n743), .Y(n440) );
  INVX1 U2691 ( .A(n735), .Y(n448) );
  INVX1 U2692 ( .A(n745), .Y(n438) );
  INVX1 U2693 ( .A(n725), .Y(n458) );
  INVX1 U2694 ( .A(n741), .Y(n442) );
  INVX1 U2695 ( .A(n721), .Y(n462) );
  INVX1 U2696 ( .A(n1066), .Y(n869) );
  INVX1 U2697 ( .A(n2346), .Y(n874) );
  INVX1 U2698 ( .A(n1072), .Y(n863) );
  INVX1 U2699 ( .A(n1068), .Y(n867) );
  INVX1 U2700 ( .A(n1070), .Y(n865) );
  INVX1 U2701 ( .A(n1069), .Y(n866) );
  INVX1 U2702 ( .A(n1071), .Y(n864) );
  INVX1 U2703 ( .A(n1073), .Y(n862) );
  INVX1 U2704 ( .A(n1067), .Y(n868) );
  INVX1 U2705 ( .A(n2401), .Y(n2395) );
  INVX1 U2706 ( .A(n2401), .Y(n2394) );
  INVX1 U2707 ( .A(n2440), .Y(n2437) );
  INVX1 U2708 ( .A(n2442), .Y(n2431) );
  INVX1 U2709 ( .A(n2420), .Y(n2413) );
  INVX1 U2710 ( .A(n2420), .Y(n2414) );
  INVX1 U2711 ( .A(n2421), .Y(n2411) );
  INVX1 U2712 ( .A(n2447), .Y(n2458) );
  INVX1 U2713 ( .A(n2447), .Y(n2459) );
  INVX1 U2714 ( .A(n2388), .Y(n2392) );
  INVX1 U2715 ( .A(n2421), .Y(n2410) );
  INVX1 U2716 ( .A(n2401), .Y(n2391) );
  INVX1 U2717 ( .A(n2481), .Y(n2469) );
  INVX1 U2718 ( .A(n2422), .Y(n2409) );
  INVX1 U2719 ( .A(n2422), .Y(n2408) );
  INVX1 U2720 ( .A(n2422), .Y(n2407) );
  INVX1 U2721 ( .A(n2466), .Y(n2448) );
  INVX1 U2722 ( .A(n2485), .Y(n2492) );
  INVX1 U2723 ( .A(n2503), .Y(n2489) );
  INVX1 U2724 ( .A(n2504), .Y(n2486) );
  INVX1 U2725 ( .A(n2400), .Y(n2399) );
  INVX1 U2726 ( .A(n2463), .Y(n2462) );
  INVX1 U2727 ( .A(n2507), .Y(n2517) );
  INVX1 U2728 ( .A(n2507), .Y(n2518) );
  INVX1 U2729 ( .A(n2525), .Y(n2516) );
  INVX1 U2730 ( .A(n2507), .Y(n2514) );
  INVX1 U2731 ( .A(n2524), .Y(n2511) );
  INVX1 U2732 ( .A(n2402), .Y(n2389) );
  INVX1 U2733 ( .A(n2423), .Y(n2440) );
  INVX1 U2734 ( .A(n2423), .Y(n2441) );
  INVX1 U2735 ( .A(n2423), .Y(n2442) );
  INVX1 U2736 ( .A(SH[7]), .Y(n2400) );
  INVX1 U2737 ( .A(SH[7]), .Y(n2401) );
  INVX1 U2738 ( .A(n2403), .Y(n2419) );
  INVX1 U2739 ( .A(n2403), .Y(n2420) );
  INVX1 U2740 ( .A(n2403), .Y(n2421) );
  INVX1 U2741 ( .A(n2445), .Y(n2463) );
  INVX1 U2742 ( .A(n2445), .Y(n2464) );
  INVX1 U2743 ( .A(n2424), .Y(n2443) );
  INVX1 U2744 ( .A(n2446), .Y(n2465) );
  INVX1 U2745 ( .A(n2404), .Y(n2422) );
  INVX1 U2746 ( .A(SH[2]), .Y(n2501) );
  INVX1 U2747 ( .A(n2424), .Y(n2444) );
  INVX1 U2748 ( .A(n2484), .Y(n2503) );
  INVX1 U2749 ( .A(n2525), .Y(n2508) );
  INVX1 U2750 ( .A(n2422), .Y(n2406) );
  INVX1 U2751 ( .A(n1424), .Y(n1239) );
  INVX1 U2752 ( .A(n1425), .Y(n1238) );
  INVX1 U2753 ( .A(n2367), .Y(n1240) );
  INVX1 U2754 ( .A(n2425), .Y(n2423) );
  INVX1 U2755 ( .A(n2405), .Y(n2403) );
  INVX1 U2756 ( .A(n2447), .Y(n2445) );
  INVX1 U2757 ( .A(n2425), .Y(n2424) );
  INVX1 U2758 ( .A(n2505), .Y(n2523) );
  INVX1 U2759 ( .A(n2447), .Y(n2446) );
  INVX1 U2760 ( .A(n2405), .Y(n2404) );
  INVX1 U2761 ( .A(n2506), .Y(n2524) );
  OR2X1 U2762 ( .A(SH[15]), .B(SH[13]), .Y(n1801) );
  INVX1 U2763 ( .A(n2485), .Y(n2484) );
  INVX1 U2764 ( .A(n2387), .Y(n2402) );
  INVX1 U2765 ( .A(n2388), .Y(n2387) );
  INVX1 U2766 ( .A(n2507), .Y(n2505) );
  INVX1 U2767 ( .A(n2507), .Y(n2506) );
  OR2X1 U2768 ( .A(SH[9]), .B(SH[8]), .Y(n1804) );
  INVX1 U2769 ( .A(A[87]), .Y(n1689) );
  INVX1 U2770 ( .A(A[112]), .Y(n1714) );
  INVX1 U2771 ( .A(A[86]), .Y(n1688) );
  INVX1 U2772 ( .A(A[117]), .Y(n1719) );
  INVX1 U2773 ( .A(A[84]), .Y(n1686) );
  INVX1 U2774 ( .A(A[34]), .Y(n1636) );
  INVX1 U2775 ( .A(A[64]), .Y(n1666) );
  INVX1 U2776 ( .A(A[16]), .Y(n1618) );
  INVX1 U2777 ( .A(A[5]), .Y(n1607) );
  INVX1 U2778 ( .A(A[4]), .Y(n1606) );
  INVX1 U2779 ( .A(A[66]), .Y(n1668) );
  INVX1 U2780 ( .A(A[88]), .Y(n1690) );
  INVX1 U2781 ( .A(A[46]), .Y(n1648) );
  INVX1 U2782 ( .A(A[114]), .Y(n1716) );
  INVX1 U2783 ( .A(A[17]), .Y(n1619) );
  INVX1 U2784 ( .A(A[36]), .Y(n1638) );
  INVX1 U2785 ( .A(A[116]), .Y(n1718) );
  INVX1 U2786 ( .A(A[133]), .Y(n1735) );
  INVX1 U2787 ( .A(A[151]), .Y(n1753) );
  INVX1 U2788 ( .A(A[131]), .Y(n1733) );
  INVX1 U2789 ( .A(A[90]), .Y(n1692) );
  INVX1 U2790 ( .A(A[167]), .Y(n1769) );
  INVX1 U2791 ( .A(A[120]), .Y(n1722) );
  INVX1 U2792 ( .A(A[54]), .Y(n1656) );
  INVX1 U2793 ( .A(A[110]), .Y(n1712) );
  INVX1 U2794 ( .A(A[111]), .Y(n1713) );
  INVX1 U2795 ( .A(A[69]), .Y(n1671) );
  INVX1 U2796 ( .A(A[118]), .Y(n1720) );
  INVX1 U2797 ( .A(A[74]), .Y(n1676) );
  INVX1 U2798 ( .A(A[3]), .Y(n1605) );
  INVX1 U2799 ( .A(A[132]), .Y(n1734) );
  INVX1 U2800 ( .A(A[150]), .Y(n1752) );
  INVX1 U2801 ( .A(A[153]), .Y(n1755) );
  INVX1 U2802 ( .A(A[161]), .Y(n1763) );
  INVX1 U2803 ( .A(A[68]), .Y(n1670) );
  INVX1 U2804 ( .A(A[125]), .Y(n1727) );
  INVX1 U2805 ( .A(A[2]), .Y(n1604) );
  INVX1 U2806 ( .A(A[152]), .Y(n1754) );
  INVX1 U2807 ( .A(A[19]), .Y(n1621) );
  INVX1 U2808 ( .A(A[163]), .Y(n1765) );
  INVX1 U2809 ( .A(A[130]), .Y(n1732) );
  INVX1 U2810 ( .A(A[166]), .Y(n1768) );
  INVX1 U2811 ( .A(A[82]), .Y(n1684) );
  INVX1 U2812 ( .A(A[98]), .Y(n1700) );
  INVX1 U2813 ( .A(A[18]), .Y(n1620) );
  INVX1 U2814 ( .A(A[28]), .Y(n1630) );
  INVX1 U2815 ( .A(A[155]), .Y(n1757) );
  INVX1 U2816 ( .A(A[149]), .Y(n1751) );
  INVX1 U2817 ( .A(A[94]), .Y(n1696) );
  INVX1 U2818 ( .A(A[40]), .Y(n1642) );
  INVX1 U2819 ( .A(A[99]), .Y(n1701) );
  INVX1 U2820 ( .A(A[100]), .Y(n1702) );
  INVX1 U2821 ( .A(A[75]), .Y(n1677) );
  INVX1 U2822 ( .A(A[169]), .Y(n1771) );
  INVX1 U2823 ( .A(A[26]), .Y(n1628) );
  INVX1 U2824 ( .A(A[122]), .Y(n1724) );
  INVX1 U2825 ( .A(A[52]), .Y(n1654) );
  INVX1 U2826 ( .A(A[24]), .Y(n1626) );
  INVX1 U2827 ( .A(A[23]), .Y(n1625) );
  INVX1 U2828 ( .A(A[22]), .Y(n1624) );
  INVX1 U2829 ( .A(A[6]), .Y(n1608) );
  INVX1 U2830 ( .A(A[96]), .Y(n1698) );
  INVX1 U2831 ( .A(A[70]), .Y(n1672) );
  INVX1 U2832 ( .A(A[72]), .Y(n1674) );
  INVX1 U2833 ( .A(A[42]), .Y(n1644) );
  INVX1 U2834 ( .A(A[39]), .Y(n1641) );
  INVX1 U2835 ( .A(A[124]), .Y(n1726) );
  INVX1 U2836 ( .A(A[56]), .Y(n1658) );
  INVX1 U2837 ( .A(A[25]), .Y(n1627) );
  INVX1 U2838 ( .A(A[7]), .Y(n1609) );
  INVX1 U2839 ( .A(A[139]), .Y(n1741) );
  INVX1 U2840 ( .A(A[157]), .Y(n1759) );
  INVX1 U2841 ( .A(A[38]), .Y(n1640) );
  INVX1 U2842 ( .A(A[168]), .Y(n1770) );
  INVX1 U2843 ( .A(A[162]), .Y(n1764) );
  INVX1 U2844 ( .A(A[154]), .Y(n1756) );
  INVX1 U2845 ( .A(A[148]), .Y(n1750) );
  INVX1 U2846 ( .A(A[123]), .Y(n1725) );
  INVX1 U2847 ( .A(A[27]), .Y(n1629) );
  INVX1 U2848 ( .A(A[140]), .Y(n1742) );
  INVX1 U2849 ( .A(A[15]), .Y(n1617) );
  INVX1 U2850 ( .A(A[20]), .Y(n1622) );
  INVX1 U2851 ( .A(A[32]), .Y(n1634) );
  INVX1 U2852 ( .A(A[14]), .Y(n1616) );
  INVX1 U2853 ( .A(A[138]), .Y(n1740) );
  INVX1 U2854 ( .A(A[141]), .Y(n1743) );
  INVX1 U2855 ( .A(A[156]), .Y(n1758) );
  INVX1 U2856 ( .A(A[57]), .Y(n1659) );
  INVX1 U2857 ( .A(A[21]), .Y(n1623) );
  INVX1 U2858 ( .A(A[33]), .Y(n1635) );
  INVX1 U2859 ( .A(A[44]), .Y(n1646) );
  INVX1 U2860 ( .A(A[1]), .Y(n1603) );
  INVX1 U2861 ( .A(A[0]), .Y(n1602) );
  INVX1 U2862 ( .A(A[45]), .Y(n1647) );
  INVX1 U2863 ( .A(A[48]), .Y(n1650) );
  INVX1 U2864 ( .A(A[143]), .Y(n1745) );
  INVX1 U2865 ( .A(A[76]), .Y(n1678) );
  INVX1 U2866 ( .A(A[108]), .Y(n1710) );
  INVX1 U2867 ( .A(A[113]), .Y(n1715) );
  INVX1 U2868 ( .A(A[115]), .Y(n1717) );
  INVX1 U2869 ( .A(A[92]), .Y(n1694) );
  INVX1 U2870 ( .A(A[67]), .Y(n1669) );
  INVX1 U2871 ( .A(A[37]), .Y(n1639) );
  INVX1 U2872 ( .A(A[65]), .Y(n1667) );
  INVX1 U2873 ( .A(A[89]), .Y(n1691) );
  INVX1 U2874 ( .A(A[35]), .Y(n1637) );
  INVX1 U2875 ( .A(A[47]), .Y(n1649) );
  INVX1 U2876 ( .A(A[105]), .Y(n1707) );
  INVX1 U2877 ( .A(A[50]), .Y(n1652) );
  INVX1 U2878 ( .A(A[85]), .Y(n1687) );
  INVX1 U2879 ( .A(A[142]), .Y(n1744) );
  INVX1 U2880 ( .A(A[58]), .Y(n1660) );
  INVX1 U2881 ( .A(A[80]), .Y(n1682) );
  INVX1 U2882 ( .A(A[104]), .Y(n1706) );
  INVX1 U2883 ( .A(A[51]), .Y(n1653) );
  INVX1 U2884 ( .A(A[91]), .Y(n1693) );
  INVX1 U2885 ( .A(A[173]), .Y(n1775) );
  INVX1 U2886 ( .A(A[55]), .Y(n1657) );
  INVX1 U2887 ( .A(A[81]), .Y(n1683) );
  INVX1 U2888 ( .A(A[119]), .Y(n1721) );
  INVX1 U2889 ( .A(A[121]), .Y(n1723) );
  INVX1 U2890 ( .A(A[158]), .Y(n1760) );
  INVX1 U2891 ( .A(A[95]), .Y(n1697) );
  INVX1 U2892 ( .A(A[83]), .Y(n1685) );
  INVX1 U2893 ( .A(A[101]), .Y(n1703) );
  INVX1 U2894 ( .A(A[41]), .Y(n1643) );
  INVX1 U2895 ( .A(A[29]), .Y(n1631) );
  INVX1 U2896 ( .A(A[159]), .Y(n1761) );
  INVX1 U2897 ( .A(A[172]), .Y(n1774) );
  INVX1 U2898 ( .A(A[71]), .Y(n1673) );
  INVX1 U2899 ( .A(A[53]), .Y(n1655) );
  INVX1 U2900 ( .A(A[97]), .Y(n1699) );
  INVX1 U2901 ( .A(A[73]), .Y(n1675) );
  INVX1 U2902 ( .A(A[43]), .Y(n1645) );
  INVX1 U2903 ( .A(A[78]), .Y(n1680) );
  INVX1 U2904 ( .A(A[145]), .Y(n1747) );
  INVX1 U2905 ( .A(A[106]), .Y(n1708) );
  INVX1 U2906 ( .A(A[49]), .Y(n1651) );
  INVX1 U2907 ( .A(A[144]), .Y(n1746) );
  INVX1 U2908 ( .A(A[77]), .Y(n1679) );
  INVX1 U2909 ( .A(A[93]), .Y(n1695) );
  INVX1 U2910 ( .A(A[109]), .Y(n1711) );
  INVX1 U2911 ( .A(A[59]), .Y(n1661) );
  INVX1 U2912 ( .A(A[107]), .Y(n1709) );
  INVX1 U2913 ( .A(A[79]), .Y(n1681) );
  INVX1 U2914 ( .A(A[63]), .Y(n1665) );
  INVX1 U2915 ( .A(A[127]), .Y(n1729) );
  INVX1 U2916 ( .A(A[60]), .Y(n1662) );
  INVX1 U2917 ( .A(A[30]), .Y(n1632) );
  INVX1 U2918 ( .A(A[12]), .Y(n1614) );
  INVX1 U2919 ( .A(A[62]), .Y(n1664) );
  INVX1 U2920 ( .A(A[102]), .Y(n1704) );
  INVX1 U2921 ( .A(A[13]), .Y(n1615) );
  INVX1 U2922 ( .A(A[135]), .Y(n1737) );
  INVX1 U2923 ( .A(A[134]), .Y(n1736) );
  INVX1 U2924 ( .A(A[10]), .Y(n1612) );
  INVX1 U2925 ( .A(A[11]), .Y(n1613) );
  INVX1 U2926 ( .A(A[137]), .Y(n1739) );
  INVX1 U2927 ( .A(A[126]), .Y(n1728) );
  INVX1 U2928 ( .A(A[175]), .Y(n1777) );
  INVX1 U2929 ( .A(A[136]), .Y(n1738) );
  INVX1 U2930 ( .A(A[8]), .Y(n1610) );
  INVX1 U2931 ( .A(A[9]), .Y(n1611) );
  INVX1 U2932 ( .A(A[146]), .Y(n1748) );
  INVX1 U2933 ( .A(A[103]), .Y(n1705) );
  INVX1 U2934 ( .A(A[31]), .Y(n1633) );
  INVX1 U2935 ( .A(A[147]), .Y(n1749) );
  INVX1 U2936 ( .A(A[61]), .Y(n1663) );
  INVX1 U2937 ( .A(A[170]), .Y(n1772) );
  INVX1 U2938 ( .A(A[128]), .Y(n1730) );
  INVX1 U2939 ( .A(A[129]), .Y(n1731) );
  INVX1 U2940 ( .A(A[165]), .Y(n1767) );
  INVX1 U2941 ( .A(A[164]), .Y(n1766) );
  INVX1 U2942 ( .A(A[160]), .Y(n1762) );
  INVX1 U2943 ( .A(A[176]), .Y(n1778) );
  INVX1 U2944 ( .A(A[177]), .Y(n1779) );
  INVX1 U2945 ( .A(A[174]), .Y(n1776) );
  INVX1 U2946 ( .A(A[171]), .Y(n1773) );
  INVX1 U2947 ( .A(A[179]), .Y(n1781) );
  INVX1 U2948 ( .A(A[178]), .Y(n1780) );
  AND2X2 U2949 ( .A(n2251), .B(n2333), .Y(B[43]) );
  AND2X2 U2950 ( .A(n2284), .B(n2381), .Y(B[31]) );
  AND2X2 U2951 ( .A(n2239), .B(n2379), .Y(B[25]) );
  AND2X2 U2952 ( .A(n2283), .B(n2318), .Y(B[29]) );
  AND2X2 U2953 ( .A(n2241), .B(n2381), .Y(B[27]) );
  AND2X2 U2954 ( .A(n2280), .B(n2315), .Y(B[22]) );
  AND2X2 U2955 ( .A(n2278), .B(n2316), .Y(B[20]) );
  AND2X2 U2956 ( .A(n2237), .B(n2382), .Y(B[16]) );
  AND2X2 U2957 ( .A(n2243), .B(n2381), .Y(B[34]) );
  AND2X2 U2958 ( .A(n2244), .B(n2333), .Y(B[35]) );
  AND2X2 U2959 ( .A(n2275), .B(n2384), .Y(B[17]) );
  AND2X2 U2960 ( .A(n2273), .B(n2379), .Y(B[14]) );
  AND2X2 U2961 ( .A(n2307), .B(n2223), .Y(B[32]) );
  AND2X2 U2962 ( .A(n2269), .B(n2380), .Y(B[6]) );
  AND2X2 U2963 ( .A(n2276), .B(n2315), .Y(B[18]) );
  AND2X2 U2964 ( .A(n2363), .B(n2380), .Y(B[0]) );
  AND2X2 U2965 ( .A(n2266), .B(n2292), .Y(n2372) );
  AND2X2 U2966 ( .A(n2377), .B(n2378), .Y(n2373) );
  AND2X2 U2967 ( .A(n2285), .B(n2383), .Y(B[33]) );
endmodule


module maze_router ( reset, start, clk, address, data_in, data_out, cs, we, D
 );
  output [7:0] address;
  input [7:0] data_in;
  output [7:0] data_out;
  input reset, start, clk;
  output cs, we, D;
  wire   n2219, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, addrLock, wS, wT, n2261, n2262, n2263, n2264,
         n2265, n2266, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3772, n3773,
         n3774, n4125, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4224, n4225, n4226, n4227, n7906, n8034,
         n8035, n8036, n8037, n8038, n8039, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n11043, n11045,
         n11047, n11049, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13799, n13800, n13801, n13802, n13803, n13804, n19662,
         n19663, n19664, n20534, n20535, n20536, n20537, n20538, n20539,
         n21313, n21314, n21315, n21316, n21317, n21318, n21322, n21323,
         n21324, n21325, n21328, n21329, n21331, n21332, n21334, n21335,
         n21337, n21338, n21340, n21341, n21343, n21344, n21346, n21347,
         n21349, n21350, n21352, n21353, n21355, n21356, n21358, n21359,
         n21361, n21362, n21364, n21365, n21367, n21368, n21370, n21371,
         n21373, n21374, n21376, n21377, n21379, n21380, n21382, n21383,
         n21385, n21386, n21388, n21389, n21391, n21392, n21394, n21395,
         n21397, n21398, n21400, n21401, n21403, n21404, n21406, n21407,
         n21409, n21410, n21412, n21413, n21415, n21416, n21418, n21419,
         n21421, n21422, n21424, n21425, n21427, n21428, n21430, n21431,
         n21433, n21434, n21436, n21437, n21439, n21440, n21442, n21443,
         n21445, n21446, n21448, n21449, n21451, n21452, n21454, n21455,
         n21457, n21458, n21460, n21461, n21463, n21464, n21466, n21468,
         n21470, n21471, n21473, n21474, n21476, n21477, n21479, n21480,
         n21482, n21483, n21485, n21486, n21488, n21489, n21491, n21492,
         n21494, n21495, n21497, n21498, n21500, n21501, n21503, n21504,
         n21506, n21507, n21509, n21510, n21512, n21513, n21515, n21516,
         n21518, n21519, n21521, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21852, n21854,
         n21858, n21860, n22053, n22054, n22055, n22056, n22058, n22059,
         n22060, n22063, n22064, n22066, n22067, n22068, n22071, n22072,
         n22074, n22075, n22076, n22079, n22080, n22082, n22083, n22084,
         n22087, n22088, n22090, n22091, n22092, n22093, n22095, n22096,
         n22098, n22099, n22100, n22101, n22103, n22104, n22105, n22106,
         n22107, n22108, n22111, n22112, n22114, n22115, n22116, n22117,
         n22119, n22120, n22121, n22123, n22124, n22125, n22127, n22128,
         n22131, n22132, n22133, n22135, n22136, n22137, n22139, n22140,
         n22141, n22143, n22144, n22147, n22148, n22149, n22151, n22152,
         n22153, n22155, n22156, n22157, n22159, n22160, n22161, n22163,
         n22164, n22165, n22167, n22168, n22171, n22172, n22173, n22175,
         n22176, n22179, n22180, n22181, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22223,
         n22224, n22225, n22226, n22227, n22228, n22231, n22232, n22233,
         n22234, n22235, n22236, n22239, n22240, n22242, n22243, n22244,
         n22247, n22248, n22249, n22251, n22252, n22253, n22255, n22256,
         n22257, n22259, n22260, n22261, n22263, n22264, n22267, n22268,
         n22269, n22271, n22272, n22275, n22276, n22277, n22279, n22280,
         n22281, n22283, n22284, n22285, n22287, n22288, n22289, n22291,
         n22292, n22293, n22295, n22296, n22297, n22299, n22300, n22301,
         n22303, n22304, n22305, n22308, n22309, n22323, n22324, n22325,
         n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
         n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341,
         n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
         n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
         n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
         n22374, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22435, n22436,
         n22438, n22439, n22441, n22442, n22444, n22445, n22447, n22448,
         n22450, n22451, n22453, n22454, n22456, n22457, n22459, n22460,
         n22462, n22463, n22465, n22466, n22468, n22469, n22471, n22472,
         n22474, n22475, n22477, n22478, n22480, n22481, n22483, n22484,
         n22486, n22487, n22489, n22490, n22492, n22493, n22495, n22496,
         n22498, n22499, n22501, n22502, n22504, n22505, n22507, n22508,
         n22510, n22511, n22513, n22514, n22516, n22517, n22519, n22520,
         n22522, n22523, n22525, n22526, n22528, n22529, n22531, n22532,
         n22534, n22535, n22537, n22538, n22540, n22541, n22543, n22544,
         n22546, n22547, n22549, n22550, n22552, n22553, n22555, n22556,
         n22558, n22559, n22561, n22562, n22564, n22565, n22567, n22568,
         n22570, n22571, n22573, n22574, n22576, n22577, n22579, n22580,
         n22582, n22583, n22585, n22586, n22588, n22589, n22591, n22592,
         n22594, n22595, n22597, n22598, n22600, n22601, n22603, n22604,
         n22606, n22607, n22609, n22610, n22612, n22613, n22615, n22616,
         n22618, n22619, n22621, n22622, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n13743, n13994, n14097, n14218, n14346, n14348,
         n14349, n14350, n14351, n14354, n14355, n14356, n14357, n14358,
         n14366, n14368, n14369, n14371, n14372, n14373, n14374, n14382,
         n14384, n14390, n14391, n14396, n14398, n14403, n14404, n14409,
         n14411, n14416, n14417, n14422, n14424, n14429, n14430, n14435,
         n14437, n14442, n14443, n14448, n14450, n14455, n14456, n14461,
         n14463, n14468, n14469, n14474, n14476, n14477, n14478, n14483,
         n14484, n14489, n14495, n14496, n14501, n14507, n14508, n14513,
         n14519, n14520, n14525, n14531, n14532, n14537, n14543, n14544,
         n14549, n14555, n14556, n14561, n14567, n14568, n14573, n14575,
         n14576, n14581, n14582, n14587, n14593, n14594, n14599, n14605,
         n14606, n14611, n14617, n14618, n14623, n14629, n14630, n14635,
         n14641, n14642, n14647, n14653, n14654, n14659, n14665, n14666,
         n14671, n14673, n14674, n14675, n14680, n14681, n14686, n14692,
         n14693, n14698, n14704, n14705, n14710, n14716, n14717, n14722,
         n14728, n14729, n14734, n14740, n14741, n14746, n14752, n14753,
         n14758, n14764, n14765, n14770, n14772, n14773, n14778, n14779,
         n14784, n14790, n14791, n14796, n14802, n14803, n14808, n14814,
         n14815, n14820, n14826, n14827, n14832, n14838, n14839, n14844,
         n14850, n14851, n14856, n14862, n14863, n14868, n14870, n14871,
         n14876, n14877, n14882, n14888, n14889, n14894, n14900, n14901,
         n14906, n14912, n14913, n14918, n14924, n14925, n14930, n14936,
         n14937, n14942, n14948, n14949, n14954, n14960, n14961, n14966,
         n14968, n14969, n14974, n14975, n14980, n14986, n14987, n14992,
         n14998, n14999, n15004, n15010, n15011, n15016, n15022, n15023,
         n15028, n15034, n15035, n15040, n15046, n15047, n15052, n15058,
         n15059, n15064, n15066, n15071, n15072, n15077, n15083, n15084,
         n15089, n15095, n15096, n15101, n15107, n15108, n15113, n15119,
         n15120, n15125, n15131, n15132, n15137, n15143, n15144, n15149,
         n15155, n15156, n15157, n15167, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15194, n15195, n15196, n15201, n15202, n15204, n15205,
         n15222, n15226, n15235, n15245, n15256, n15260, n15269, n15279,
         n15283, n15293, n15302, n15306, n15316, n15325, n15329, n15339,
         n15348, n15352, n15362, n15373, n15377, n15387, n15397, n15401,
         n15411, n15420, n15424, n15434, n15442, n15446, n15456, n15464,
         n15469, n15478, n15486, n15490, n15500, n15508, n15512, n15521,
         n15529, n15535, n15544, n15552, n15566, n15574, n15580, n15589,
         n15597, n15601, n15611, n15618, n15623, n15632, n15639, n15644,
         n15653, n15660, n15665, n15674, n15681, n15686, n15695, n15702,
         n15707, n15716, n15724, n15729, n15738, n15746, n15751, n15760,
         n15767, n15772, n15781, n15788, n15793, n15802, n15809, n15814,
         n15823, n15830, n15835, n15844, n15851, n15856, n15865, n15872,
         n15873, n15879, n15880, n15887, n15897, n15899, n15900, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15955, n15956, n15957, n15958, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15970, n15971,
         n15972, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15985, n15986, n15987, n15988, n15989, n15992, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16017, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16030, n16031, n16032, n16034, n16035, n16036, n16039, n16044,
         n16051, n16052, n16053, n16055, n16056, n16057, n16059, n16060,
         n16061, n16062, n16063, n16066, n16071, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16106, n16107, n16108, n16109, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16121, n16122, n16123,
         n16128, n16129, n16130, n16132, n16133, n16134, n16136, n16137,
         n16138, n16139, n16140, n16143, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16175, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16187, n16188, n16189,
         n16190, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16202, n16203, n16204, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16217, n16218, n16219, n16220, n16221, n16224,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16242, n16243, n16244, n16245, n16247, n16269, n16280, n16281,
         net53176, net53596, net53601, net53623, net53785, net64168, net89744,
         net89759, net89777, net89785, net89806, net90010, net90052, net90053,
         net90054, net90055, net90071, net94645, net94647, net94649, net95105,
         net95147, net95156, net95303, net95456, net95457, net95464, net95480,
         net96340, net96604, net96600, net96598, net96596, net96592, net96588,
         net96586, net96584, net96582, net96578, net96576, net96574, net96572,
         net96570, net96568, net96566, net96564, net96562, net96560, net96558,
         alt5_net95652, alt5_net95654, alt5_net95656, alt5_net95658,
         alt5_net95662, alt5_net95664, alt5_net95666, alt5_net95668,
         alt5_net95670, alt5_net95676, alt14_net96326, alt14_net96328,
         alt14_net96302, alt14_net96304, alt14_net96306, alt14_net96296,
         alt14_net96264, alt14_net96268, alt14_net96230, alt14_net96236,
         alt14_net96238, alt14_net96248, alt14_net96250, alt14_net96258,
         alt14_net55935, alt14_net55927, alt14_net55921, alt14_net6254,
         alt14_net6253, alt14_net6192, alt14_net6191, alt14_net6130,
         alt14_net6129, alt14_net6006, alt14_net6005, net102091, net103671,
         net103869, net104480, net104479, net104600, net105779, net105778,
         net105788, net105787, net105786, net105822, net105821, net105819,
         net105816, net105815, net105814, net105813, net105810, net105808,
         net105807, net105803, net105802, net105801, net105800, net105799,
         net105798, net105797, net105796, net105795, net105794, net105793,
         net105859, net105857, net106018, net106017, net107094, net107091,
         net107090, net107088, net107082, net107078, net107076, net107074,
         net107063, net107061, net108311, net108471, net108478, net108619,
         net108653, net108805, net108804, net108803, net109176, net109385,
         net109417, net109440, net109469, net109485, net109512, net109585,
         net109766, net109824, net110246, net110320, net110411, net110410,
         net110421, net110687, net110686, net110685, net110809, net110815,
         net110814, net110825, net110927, net110926, net111205, net111222,
         net111237, net111332, net111600, net111628, net111984, net112181,
         net112188, net112192, net112194, net112202, net112859, net112858,
         net113308, net113321, net113687, net113686, net113955, net113954,
         net114151, net114244, net114253, net114252, net114546, net114723,
         net114744, net114808, net114916, net115535, net115619, net115636,
         net115635, net116755, net116754, net116760, net116777, net116776,
         net116925, net116949, net117076, net117217, net117301, net124030,
         net124029, net125067, net125066, net137490, net137489, net137830,
         net138161, net138174, net142478, net142728, net142789, net142788,
         net143010, net143109, net144199, net145105, net145121, net145295,
         net146640, net146826, net146838, net147379, net147507, net147506,
         net147505, net147504, net147502, net147501, net147500, net147499,
         net147498, net147497, net147496, net147495, net147494, net147493,
         net147492, net147490, net147481, net147761, net147983, net149749,
         net149764, net149842, net149850, net149863, net149862, net149877,
         net149876, net149909, net149922, net149936, net149941, net149940,
         net149947, net149983, net149982, net149986, net150046, net150085,
         net150126, net150130, net150133, net150132, net150220, net150245,
         net150251, net150253, net150331, net150330, net150376, net150385,
         net150650, net150787, net151212, net151429, net151617, net151626,
         net151629, net151633, net151632, net151649, net151652, net151662,
         net151697, net151696, net151710, net151709, net151738, net151741,
         net151751, net151801, net151812, net151814, net151834, net151833,
         net151840, net151875, net151887, net151886, net151977, net147735,
         n21834, net90056, net150261, net142746, n4223, net95477, net90064,
         net143040, net139028, net105988, n14360, n14359, alt14_net96276,
         net95482, net143105, n4126, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21319, n21320,
         n21321, n21326, n21327, n21330, n21333, n21336, n21339, n21342,
         n21345, n21348, n21351, n21354, n21357, n21360, n21363, n21366,
         n21369, n21372, n21375, n21378, n21381, n21384, n21387, n21390,
         n21393, n21396, n21399, n21402, n21405, n21408, n21411, n21414,
         n21417, n21420, n21423, n21426, n21429, n21432, n21435, n21438,
         n21441, n21444, n21447, n21450, n21453, n21456, n21459, n21462,
         n21465, n21467, n21469, n21472, n21475, n21478, n21481, n21484,
         n21487, n21490, n21493, n21496, n21499, n21502, n21505, n21508,
         n21511, n21514, n21517, n21520, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21666, n21699, n21767, n21782, n21801, n21848, n21849,
         n21850, n21851, n21853, n21855, n21856, n21857, n21859, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22057,
         n22061, n22062, n22065, n22069, n22070, n22073, n22077, n22078,
         n22081, n22085, n22086, n22089, n22094, n22097, n22102, n22109,
         n22110, n22113, n22118, n22122, n22126, n22129, n22130, n22134,
         n22138, n22142, n22145, n22146, n22150, n22154, n22158, n22162,
         n22166, n22169, n22170, n22174, n22177, n22178, n22182, n22190,
         n22198, n22206, n22214, n22222, n22229, n22230, n22237, n22238,
         n22241, n22245, n22246, n22250, n22254, n22258, n22262, n22265,
         n22266, n22270, n22273, n22274, n22278, n22282, n22286, n22290,
         n22294, n22298, n22302, n22306, n22307, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22375, n22420, n22421, n22422, n22423, n22424,
         n22434, n22437, n22440, n22443, n22446, n22449, n22452, n22455,
         n22458, n22461, n22464, n22467, n22470, n22473, n22476, n22479,
         n22482, n22485, n22488, n22491, n22494, n22497, n22500, n22503,
         n22506, n22509, n22512, n22515, n22518, n22521, n22524, n22527,
         n22530, n22533, n22536, n22539, n22542, n22545, n22548, n22551,
         n22554, n22557, n22560, n22563, n22566, n22569, n22572, n22575,
         n22578, n22581, n22584, n22587, n22590, n22593, n22596, n22599,
         n22602, n22605, n22608, n22611, n22614, n22617, n22620, n22623,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
         n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
         n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
         n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773,
         n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
         n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
         n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
         n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
         n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
         n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
         n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
         n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
         n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845,
         n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
         n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
         n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
         n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
         n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
         n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
         n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
         n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
         n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917,
         n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
         n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
         n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
         n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
         n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
         n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
         n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
         n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
         n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
         n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
         n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
         n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
         n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
         n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
         n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
         n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101,
         n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109,
         n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
         n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
         n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
         n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181,
         n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
         n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
         n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205,
         n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
         n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
         n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
         n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
         n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
         n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
         n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
         n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
         n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
         n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
         n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
         n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301,
         n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
         n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
         n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
         n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
         n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
         n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
         n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
         n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
         n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373,
         n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
         n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
         n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
         n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
         n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
         n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
         n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
         n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
         n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
         n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
         n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
         n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
         n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
         n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
         n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
         n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
         n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
         n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
         n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
         n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
         n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
         n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
         n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
         n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
         n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
         n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
         n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
         n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
         n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
         n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
         n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
         n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
         n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
         n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
         n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
         n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
         n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
         n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
         n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
         n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
         n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
         n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
         n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
         n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
         n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
         n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
         n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
         n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
         n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
         n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
         n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
         n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
         n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
         n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
         n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
         n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165,
         n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
         n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
         n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
         n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
         n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
         n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
         n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
         n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
         n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237,
         n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
         n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
         n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
         n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
         n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
         n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
         n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
         n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
         n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309,
         n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
         n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
         n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
         n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
         n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
         n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357,
         n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
         n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
         n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381,
         n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
         n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
         n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405,
         n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
         n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
         n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429,
         n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
         n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
         n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
         n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
         n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
         n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
         n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
         n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
         n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
         n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
         n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
         n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
         n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573,
         n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
         n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
         n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
         n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
         n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
         n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621,
         n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
         n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
         n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
         n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
         n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
         n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
         n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
         n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
         n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
         n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
         n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
         n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717,
         n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725,
         n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
         n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
         n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
         n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
         n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
         n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
         n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797,
         n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
         n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
         n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
         n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
         n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837,
         n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
         n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
         n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861,
         n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869,
         n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
         n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
         n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
         n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
         n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909,
         n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
         n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
         n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933,
         n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941,
         n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
         n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
         n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
         n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
         n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981,
         n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
         n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
         n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005,
         n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
         n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
         n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
         n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
         n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
         n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053,
         n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
         n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
         n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
         n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
         n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
         n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
         n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197,
         n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
         n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
         n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
         n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
         n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
         n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
         n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
         n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
         n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
         n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301,
         n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
         n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
         n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
         n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
         n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341,
         n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
         n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
         n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
         n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
         n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
         n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
         n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413,
         n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
         n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
         n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
         n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445,
         n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
         n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
         n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
         n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
         n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485,
         n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
         n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
         n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
         n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517,
         n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
         n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
         n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
         n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549,
         n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557,
         n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
         n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
         n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581,
         n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589,
         n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
         n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
         n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
         n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621,
         n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629,
         n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
         n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661,
         n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
         n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677,
         n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
         n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693,
         n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701,
         n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
         n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
         n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725,
         n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733,
         n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
         n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749,
         n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
         n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
         n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773,
         n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
         n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
         n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
         n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
         n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
         n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821,
         n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
         n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
         n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
         n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
         n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
         n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
         n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893,
         n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
         n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925,
         n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
         n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
         n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
         n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
         n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965,
         n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
         n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
         n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
         n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013,
         n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
         n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
         n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
         n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
         n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
         n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133,
         n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
         n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
         n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165,
         n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
         n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
         n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
         n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237,
         n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277,
         n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
         n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
         n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309,
         n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
         n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
         n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
         n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349,
         n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
         n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
         n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
         n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
         n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397,
         n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
         n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
         n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421,
         n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
         n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
         n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445,
         n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453,
         n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
         n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469,
         n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
         n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
         n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493,
         n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501,
         n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
         n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
         n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
         n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
         n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541,
         n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
         n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
         n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
         n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589,
         n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
         n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
         n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
         n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
         n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
         n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
         n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
         n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
         n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
         n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
         n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
         n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117,
         n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
         n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
         n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
         n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
         n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
         n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
         n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
         n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
         n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
         n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
         n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
         n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
         n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
         n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
         n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
         n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
         n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381,
         n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389,
         n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
         n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421,
         n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
         n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
         n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445,
         n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453,
         n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461,
         n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
         n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
         n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
         n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
         n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501,
         n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
         n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
         n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
         n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
         n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
         n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
         n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597,
         n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
         n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
         n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
         n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
         n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
         n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
         n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
         n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
         n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813,
         n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821,
         n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
         n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
         n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
         n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
         n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
         n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
         n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
         n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
         n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
         n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
         n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037,
         n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
         n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
         n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
         n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
         n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
         n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109,
         n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
         n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
         n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
         n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
         n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
         n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
         n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
         n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
         n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389,
         n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
         n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
         n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
         n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437,
         n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445,
         n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469,
         n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
         n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
         n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
         n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
         n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509,
         n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517,
         n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
         n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533,
         n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541,
         n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
         n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
         n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
         n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581,
         n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
         n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
         n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
         n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
         n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
         n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653,
         n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
         n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669,
         n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677,
         n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685,
         n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
         n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
         n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
         n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717,
         n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725,
         n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733,
         n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741,
         n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749,
         n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757,
         n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
         n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773,
         n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
         n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789,
         n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797,
         n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805,
         n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813,
         n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821,
         n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829,
         n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837,
         n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845,
         n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
         n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861,
         n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869,
         n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877,
         n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885,
         n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893,
         n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901,
         n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909,
         n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
         n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
         n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933,
         n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941,
         n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949,
         n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957,
         n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965,
         n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973,
         n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981,
         n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
         n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997,
         n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005,
         n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013,
         n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021,
         n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029,
         n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037,
         n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045,
         n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
         n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061,
         n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069,
         n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
         n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085,
         n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
         n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
         n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109,
         n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117,
         n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
         n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
         n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
         n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149,
         n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157,
         n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
         n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173,
         n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181,
         n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189,
         n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
         n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205,
         n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213,
         n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221,
         n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229,
         n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237,
         n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245,
         n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253,
         n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261,
         n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
         n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277,
         n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
         n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293,
         n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301,
         n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309,
         n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317,
         n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325,
         n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333,
         n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
         n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349,
         n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357,
         n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365,
         n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373,
         n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381,
         n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389,
         n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397,
         n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405,
         n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
         n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
         n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
         n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
         n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
         n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453,
         n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461,
         n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469,
         n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
         n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
         n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493,
         n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501,
         n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509,
         n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517,
         n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525,
         n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533,
         n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541,
         n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549,
         n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
         n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565,
         n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573,
         n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581,
         n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589,
         n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597,
         n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605,
         n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613,
         n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621,
         n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
         n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637,
         n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645,
         n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653,
         n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661,
         n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669,
         n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677,
         n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685,
         n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693,
         n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
         n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709,
         n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
         n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
         n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733,
         n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
         n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749,
         n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757,
         n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765,
         n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
         n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781,
         n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
         n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797,
         n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805,
         n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813,
         n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821,
         n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829,
         n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837,
         n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
         n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853,
         n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861,
         n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869,
         n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877,
         n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885,
         n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893,
         n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901,
         n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909,
         n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
         n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925,
         n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933,
         n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941,
         n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949,
         n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957,
         n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965,
         n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973,
         n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981,
         n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989,
         n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997,
         n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005,
         n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013,
         n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021,
         n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029,
         n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037,
         n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045,
         n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053,
         n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
         n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069,
         n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077,
         n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085,
         n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093,
         n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101,
         n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109,
         n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117,
         n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125,
         n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
         n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141,
         n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
         n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157,
         n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165,
         n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173,
         n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181,
         n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189,
         n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197,
         n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
         n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213,
         n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221,
         n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229,
         n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237,
         n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
         n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253,
         n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261,
         n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269,
         n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
         n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285,
         n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
         n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301,
         n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309,
         n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317,
         n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
         n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333,
         n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341,
         n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
         n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357,
         n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365,
         n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
         n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381,
         n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389,
         n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397,
         n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405,
         n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413,
         n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
         n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429,
         n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437,
         n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445,
         n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453,
         n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461,
         n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469,
         n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477,
         n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485,
         n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
         n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501,
         n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509,
         n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517,
         n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525,
         n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533,
         n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541,
         n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549,
         n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557,
         n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
         n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573,
         n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581,
         n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589,
         n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597,
         n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605,
         n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613,
         n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621,
         n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629,
         n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
         n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645,
         n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653,
         n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661,
         n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669,
         n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677,
         n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685,
         n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693,
         n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701,
         n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709,
         n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717,
         n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725,
         n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733,
         n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741,
         n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749,
         n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757,
         n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765,
         n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773,
         n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
         n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789,
         n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797,
         n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805,
         n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813,
         n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821,
         n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829,
         n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837,
         n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845,
         n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853,
         n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861,
         n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869,
         n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877,
         n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885,
         n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893,
         n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901,
         n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909,
         n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917,
         n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925,
         n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933,
         n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941,
         n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949,
         n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957,
         n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965,
         n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973,
         n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981,
         n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989,
         n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
         n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005,
         n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013,
         n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021,
         n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029,
         n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037,
         n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
         n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053,
         n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061,
         n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069,
         n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077,
         n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085,
         n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093,
         n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101,
         n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109,
         n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117,
         n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125,
         n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133,
         n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141,
         n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149,
         n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157,
         n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165,
         n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173,
         n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181,
         n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189,
         n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197,
         n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205,
         n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213,
         n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221,
         n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229,
         n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237,
         n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245,
         n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253,
         n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261,
         n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269,
         n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277,
         n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285,
         n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293,
         n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301,
         n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309,
         n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317,
         n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325,
         n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333,
         n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341,
         n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349,
         n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357,
         n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365,
         n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373,
         n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381,
         n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389,
         n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397,
         n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405,
         n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413,
         n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421,
         n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
         n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437,
         n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445,
         n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453,
         n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461,
         n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469,
         n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
         n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485,
         n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493,
         n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501,
         n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509,
         n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517,
         n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525,
         n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533,
         n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541,
         n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549,
         n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557,
         n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565,
         n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573,
         n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581,
         n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589,
         n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597,
         n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605,
         n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613,
         n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621,
         n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629,
         n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637,
         n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
         n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653,
         n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661,
         n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669,
         n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677,
         n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685,
         n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693,
         n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701,
         n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709,
         n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717,
         n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725,
         n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733,
         n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741,
         n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749,
         n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757,
         n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765,
         n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773,
         n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781,
         n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789,
         n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797,
         n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805,
         n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813,
         n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821,
         n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829,
         n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837,
         n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845,
         n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853,
         n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861,
         n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869,
         n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877,
         n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885,
         n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893,
         n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901,
         n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909,
         n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917,
         n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925,
         n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933,
         n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941,
         n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949,
         n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957,
         n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965,
         n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973,
         n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981,
         n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989,
         n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997,
         n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005,
         n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013,
         n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021,
         n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029,
         n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037,
         n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045,
         n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053,
         n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061,
         n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069,
         n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077,
         n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085,
         n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
         n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101,
         n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109,
         n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117,
         n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125,
         n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133,
         n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141,
         n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149,
         n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157,
         n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165,
         n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173,
         n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181,
         n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189,
         n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197,
         n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205,
         n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213,
         n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221,
         n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229,
         n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237,
         n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245,
         n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253,
         n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261,
         n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269,
         n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277,
         n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285,
         n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293,
         n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301,
         n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309,
         n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317,
         n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325,
         n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333,
         n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341,
         n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349,
         n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357,
         n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
         n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373,
         n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381,
         n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389,
         n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397,
         n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405,
         n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413,
         n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421,
         n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429,
         n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437,
         n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445,
         n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453,
         n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461,
         n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469,
         n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477,
         n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485,
         n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493,
         n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501,
         n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509,
         n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517,
         n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525,
         n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533,
         n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541,
         n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549,
         n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557,
         n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565,
         n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573,
         n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581,
         n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589,
         n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597,
         n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605,
         n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613,
         n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621,
         n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629,
         n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637,
         n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
         n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
         n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661,
         n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669,
         n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677,
         n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685,
         n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693,
         n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701,
         n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709,
         n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717,
         n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725,
         n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733,
         n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
         n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749,
         n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757,
         n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765,
         n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773,
         n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781,
         n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789,
         n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797,
         n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805,
         n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813,
         n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821,
         n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829,
         n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837,
         n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845,
         n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853,
         n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861,
         n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869,
         n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877,
         n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885,
         n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893,
         n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901,
         n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909,
         n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917,
         n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925,
         n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933,
         n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941,
         n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949,
         n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957,
         n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965,
         n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973,
         n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981,
         n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989,
         n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997,
         n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005,
         n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013,
         n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021,
         n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029,
         n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037,
         n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045,
         n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053,
         n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061,
         n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069,
         n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077,
         n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085,
         n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093,
         n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101,
         n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109,
         n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117,
         n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125,
         n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133,
         n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141,
         n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149,
         n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157,
         n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165,
         n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173,
         n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181,
         n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189,
         n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197,
         n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205,
         n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213,
         n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221,
         n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229,
         n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237,
         n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245,
         n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253,
         n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261,
         n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269,
         n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277,
         n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285,
         n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293,
         n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
         n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309,
         n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317,
         n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325,
         n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333,
         n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341,
         n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349,
         n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357,
         n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365,
         n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373,
         n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381,
         n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389,
         n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397,
         n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405,
         n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
         n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421,
         n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429,
         n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437,
         n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445,
         n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453,
         n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
         n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469,
         n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477,
         n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485,
         n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493,
         n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501,
         n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509,
         n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
         n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525,
         n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
         n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541,
         n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549,
         n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557,
         n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565,
         n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573,
         n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581,
         n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
         n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597,
         n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605,
         n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613,
         n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621,
         n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
         n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637,
         n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645,
         n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653,
         n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661,
         n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669,
         n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677,
         n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685,
         n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693,
         n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701,
         n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709,
         n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717,
         n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725,
         n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733,
         n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741,
         n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749,
         n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757,
         n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765,
         n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773,
         n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781,
         n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789,
         n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797,
         n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805,
         n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813,
         n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821,
         n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829,
         n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837,
         n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845,
         n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853,
         n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861,
         n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869,
         n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877,
         n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885,
         n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893,
         n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901,
         n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909,
         n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917,
         n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925,
         n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933,
         n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941,
         n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949,
         n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957,
         n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965,
         n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973,
         n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981,
         n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989,
         n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997,
         n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005,
         n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013,
         n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021,
         n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029,
         n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037,
         n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045,
         n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053,
         n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061,
         n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069,
         n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077,
         n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085,
         n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093,
         n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101,
         n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109,
         n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117,
         n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125,
         n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133,
         n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141,
         n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149,
         n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157,
         n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165,
         n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173,
         n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181,
         n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189,
         n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197,
         n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205,
         n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213,
         n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221,
         n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229,
         n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237,
         n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245,
         n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253,
         n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261,
         n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269,
         n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277,
         n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285,
         n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293,
         n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301,
         n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309,
         n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317,
         n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325,
         n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333,
         n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341,
         n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349,
         n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357,
         n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365,
         n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373,
         n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381,
         n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389,
         n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397,
         n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405,
         n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413,
         n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
         n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429,
         n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437,
         n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445,
         n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453,
         n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461,
         n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469,
         n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477,
         n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485,
         n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493,
         n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501,
         n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509,
         n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517,
         n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525,
         n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533,
         n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541,
         n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549,
         n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557,
         n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565,
         n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573,
         n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581,
         n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589,
         n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597,
         n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605,
         n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613,
         n34614, n34615, n34616, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5;
  wire   [1:0] states;
  wire   [1:0] Setup;
  wire   [179:174] RO;
  wire   [31:0] oc;
  wire   [3:0] locTrig;
  wire   [3:0] pLoc;
  wire   [179:174] RN;
  wire   [31:0] nc;
  wire   [2:0] direct;
  wire   [5:0] S;
  wire   [383:0] grid;
  wire   [5:0] T;
  wire   [2:0] direction_line;
  wire   [2:0] direction_lee;
  wire   [5:0] loc_s2;
  wire   [2:0] invdirect_s2;
  assign address[6] = 1'b0;
  assign data_out[7] = 1'b0;
  assign data_out[6] = 1'b0;
  assign data_out[5] = 1'b0;
  assign data_out[4] = 1'b0;
  assign data_out[3] = 1'b0;
  assign data_out[2] = 1'b0;
  assign data_out[1] = 1'b0;
  assign data_out[0] = 1'b0;

  LATCH T_reg_0_ ( .CLK(n22627), .D(data_in[0]), .Q(T[0]) );
  LATCH pLoc_reg_0_ ( .CLK(n22628), .D(n11043), .Q(pLoc[0]) );
  LATCH direction_lee_reg_2_ ( .CLK(n22636), .D(n34612), .Q(direction_lee[2])
         );
  LATCH nc_reg_0_ ( .CLK(n22425), .D(n21783), .Q(nc[0]) );
  LATCH nc_reg_31_ ( .CLK(n22425), .D(n21815), .Q(nc[31]) );
  LATCH oc_reg_31_ ( .CLK(n22426), .D(n23632), .Q(oc[31]) );
  LATCH RO_reg_179_ ( .CLK(n22419), .D(n34494), .Q(RO[179]) );
  LATCH pLoc_reg_3_ ( .CLK(n22631), .D(n21240), .Q(pLoc[3]) );
  LATCH direction_line_reg_2_ ( .CLK(n22633), .D(net149842), .Q(
        direction_line[2]) );
  LATCH locTrig_reg_2_ ( .CLK(n22432), .D(n21858), .Q(locTrig[2]) );
  LATCH oc_reg_30_ ( .CLK(n22426), .D(n21846), .Q(oc[30]) );
  LATCH RO_reg_178_ ( .CLK(n22419), .D(n34493), .Q(RO[178]) );
  LATCH pLoc_reg_2_ ( .CLK(n22630), .D(n21241), .Q(pLoc[2]) );
  LATCH locTrig_reg_0_ ( .CLK(n22430), .D(n21354), .Q(locTrig[0]) );
  LATCH RN_reg_179_ ( .CLK(n22425), .D(n26598), .Q(RN[179]) );
  LATCH RO_reg_177_ ( .CLK(n22418), .D(n34460), .Q(RO[177]) );
  LATCH location_reg_3_ ( .CLK(n22632), .D(n23631), .Q(n2254) );
  LATCH RO_reg_1_ ( .CLK(n22329), .D(n21329), .Q(n3103) );
  LATCH location_reg_5_ ( .CLK(n22632), .D(n23630), .Q(n2256) );
  LATCH direct_reg_0_ ( .CLK(n22634), .D(net149941), .Q(direct[0]) );
  LATCH direct_reg_2_ ( .CLK(n22634), .D(n4125), .Q(direct[2]) );
  LATCH direction_line_reg_0_ ( .CLK(n22633), .D(net138174), .Q(
        direction_line[0]) );
  LATCH direction_line_reg_1_ ( .CLK(n22633), .D(net145121), .Q(
        direction_line[1]) );
  LATCH direct_reg_1_ ( .CLK(n22634), .D(net115619), .Q(direct[1]) );
  LATCH RO_reg_0_ ( .CLK(n22329), .D(n21328), .Q(n3102) );
  LATCH location_reg_2_ ( .CLK(n22632), .D(n21351), .Q(n2253) );
  LATCH location_reg_4_ ( .CLK(n22632), .D(n21348), .Q(n2255) );
  LATCH states_reg_1_ ( .CLK(n22327), .D(n21323), .Q(states[1]) );
  LATCH states_reg_0_ ( .CLK(n22327), .D(n21239), .Q(states[0]) );
  LATCH nc_reg_30_ ( .CLK(n22425), .D(n21814), .Q(nc[30]) );
  LATCH nc_reg_29_ ( .CLK(n22425), .D(n21813), .Q(nc[29]) );
  LATCH nc_reg_28_ ( .CLK(n22425), .D(n21812), .Q(nc[28]) );
  LATCH nc_reg_27_ ( .CLK(n22425), .D(n21811), .Q(nc[27]) );
  LATCH nc_reg_26_ ( .CLK(n22425), .D(n21810), .Q(nc[26]) );
  LATCH nc_reg_25_ ( .CLK(n22425), .D(n21809), .Q(nc[25]) );
  LATCH nc_reg_24_ ( .CLK(n22425), .D(n21808), .Q(nc[24]) );
  LATCH nc_reg_23_ ( .CLK(n22425), .D(n21807), .Q(nc[23]) );
  LATCH nc_reg_22_ ( .CLK(n22425), .D(n21806), .Q(nc[22]) );
  LATCH nc_reg_21_ ( .CLK(n22425), .D(n21805), .Q(nc[21]) );
  LATCH nc_reg_20_ ( .CLK(n22425), .D(n21804), .Q(nc[20]) );
  LATCH nc_reg_19_ ( .CLK(n22425), .D(n21803), .Q(nc[19]) );
  LATCH nc_reg_18_ ( .CLK(n22425), .D(n21802), .Q(nc[18]) );
  LATCH nc_reg_17_ ( .CLK(n22425), .D(n21800), .Q(nc[17]) );
  LATCH nc_reg_16_ ( .CLK(n22425), .D(n21799), .Q(nc[16]) );
  LATCH nc_reg_15_ ( .CLK(n22425), .D(n21798), .Q(nc[15]) );
  LATCH nc_reg_14_ ( .CLK(n22425), .D(n21797), .Q(nc[14]) );
  LATCH nc_reg_13_ ( .CLK(n22425), .D(n21796), .Q(nc[13]) );
  LATCH nc_reg_12_ ( .CLK(n22425), .D(n21795), .Q(nc[12]) );
  LATCH nc_reg_11_ ( .CLK(n22425), .D(n21794), .Q(nc[11]) );
  LATCH nc_reg_10_ ( .CLK(n22425), .D(n21793), .Q(nc[10]) );
  LATCH nc_reg_9_ ( .CLK(n22425), .D(n21792), .Q(nc[9]) );
  LATCH nc_reg_8_ ( .CLK(n22425), .D(n21791), .Q(nc[8]) );
  LATCH nc_reg_7_ ( .CLK(n22425), .D(n21790), .Q(nc[7]) );
  LATCH nc_reg_6_ ( .CLK(n22425), .D(n21789), .Q(nc[6]) );
  LATCH nc_reg_5_ ( .CLK(n22425), .D(n21788), .Q(nc[5]) );
  LATCH nc_reg_4_ ( .CLK(n22425), .D(n21787), .Q(nc[4]) );
  LATCH nc_reg_3_ ( .CLK(n22425), .D(n21786), .Q(nc[3]) );
  LATCH nc_reg_2_ ( .CLK(n22425), .D(n21785), .Q(nc[2]) );
  LATCH nc_reg_1_ ( .CLK(n22425), .D(n21784), .Q(nc[1]) );
  LATCH RN_reg_178_ ( .CLK(n22425), .D(n26624), .Q(RN[178]) );
  LATCH RN_reg_177_ ( .CLK(n22425), .D(n26650), .Q(RN[177]) );
  LATCH RN_reg_176_ ( .CLK(n22425), .D(n26682), .Q(RN[176]) );
  LATCH RN_reg_175_ ( .CLK(n22425), .D(n26717), .Q(RN[175]) );
  LATCH RN_reg_174_ ( .CLK(n22425), .D(n26766), .Q(RN[174]) );
  LATCH RN_reg_173_ ( .CLK(n22425), .D(n26823), .Q(n8229) );
  LATCH RN_reg_172_ ( .CLK(n22425), .D(n26881), .Q(n8228) );
  LATCH RN_reg_171_ ( .CLK(n22425), .D(n26950), .Q(n8227) );
  LATCH RN_reg_170_ ( .CLK(n22425), .D(n27028), .Q(n8226) );
  LATCH RN_reg_169_ ( .CLK(n22425), .D(n27123), .Q(n8225) );
  LATCH RN_reg_168_ ( .CLK(n22425), .D(n23629), .Q(n8224) );
  LATCH RN_reg_167_ ( .CLK(n22425), .D(n26580), .Q(n8223) );
  LATCH RN_reg_166_ ( .CLK(n22425), .D(n26602), .Q(n8222) );
  LATCH RN_reg_165_ ( .CLK(n22425), .D(n26628), .Q(n8221) );
  LATCH RN_reg_164_ ( .CLK(n22425), .D(n26654), .Q(n8220) );
  LATCH RN_reg_163_ ( .CLK(n22425), .D(n26686), .Q(n8219) );
  LATCH RN_reg_162_ ( .CLK(n22425), .D(n26721), .Q(n8218) );
  LATCH RN_reg_161_ ( .CLK(n22425), .D(n26770), .Q(n8217) );
  LATCH RN_reg_160_ ( .CLK(n22425), .D(n26827), .Q(n8216) );
  LATCH RN_reg_159_ ( .CLK(n22425), .D(n26885), .Q(n8215) );
  LATCH RN_reg_158_ ( .CLK(n22425), .D(n26954), .Q(n8214) );
  LATCH RN_reg_157_ ( .CLK(n22425), .D(n27032), .Q(n8213) );
  LATCH RN_reg_156_ ( .CLK(n22425), .D(n27127), .Q(n8212) );
  LATCH RN_reg_155_ ( .CLK(n22425), .D(n21345), .Q(n8211) );
  LATCH RN_reg_154_ ( .CLK(n22425), .D(n26581), .Q(n8210) );
  LATCH RN_reg_153_ ( .CLK(n22425), .D(n26603), .Q(n8209) );
  LATCH RN_reg_152_ ( .CLK(n22425), .D(n26629), .Q(n8208) );
  LATCH RN_reg_151_ ( .CLK(n22425), .D(n26655), .Q(n8207) );
  LATCH RN_reg_150_ ( .CLK(n22425), .D(n26687), .Q(n8206) );
  LATCH RN_reg_149_ ( .CLK(n22425), .D(n26722), .Q(n8205) );
  LATCH RN_reg_148_ ( .CLK(n22425), .D(n26771), .Q(n8204) );
  LATCH RN_reg_147_ ( .CLK(n22425), .D(n26828), .Q(n8203) );
  LATCH RN_reg_146_ ( .CLK(n22425), .D(n26886), .Q(n8202) );
  LATCH RN_reg_145_ ( .CLK(n22425), .D(n26955), .Q(n8201) );
  LATCH RN_reg_144_ ( .CLK(n22425), .D(n27033), .Q(n8200) );
  LATCH RN_reg_143_ ( .CLK(n22425), .D(n27128), .Q(n8199) );
  LATCH RN_reg_142_ ( .CLK(n22425), .D(n21342), .Q(n8198) );
  LATCH RN_reg_141_ ( .CLK(n22425), .D(n26577), .Q(n8197) );
  LATCH RN_reg_140_ ( .CLK(n22425), .D(n26599), .Q(n8196) );
  LATCH RN_reg_139_ ( .CLK(n22425), .D(n26625), .Q(n8195) );
  LATCH RN_reg_138_ ( .CLK(n22425), .D(n26651), .Q(n8194) );
  LATCH RN_reg_137_ ( .CLK(n22425), .D(n26683), .Q(n8193) );
  LATCH RN_reg_136_ ( .CLK(n22425), .D(n26718), .Q(n8192) );
  LATCH RN_reg_135_ ( .CLK(n22425), .D(n26767), .Q(n8191) );
  LATCH RN_reg_134_ ( .CLK(n22425), .D(n26824), .Q(n8190) );
  LATCH RN_reg_133_ ( .CLK(n22425), .D(n26882), .Q(n8189) );
  LATCH RN_reg_132_ ( .CLK(n22425), .D(n26951), .Q(n8188) );
  LATCH RN_reg_131_ ( .CLK(n22425), .D(n27029), .Q(n8187) );
  LATCH RN_reg_130_ ( .CLK(n22425), .D(n27124), .Q(n8186) );
  LATCH RN_reg_129_ ( .CLK(n22425), .D(n21339), .Q(n8185) );
  LATCH RN_reg_128_ ( .CLK(n22425), .D(n26578), .Q(n8184) );
  LATCH RN_reg_127_ ( .CLK(n22425), .D(n26600), .Q(n8183) );
  LATCH RN_reg_126_ ( .CLK(n22425), .D(n26626), .Q(n8182) );
  LATCH RN_reg_125_ ( .CLK(n22425), .D(n26652), .Q(n8181) );
  LATCH RN_reg_124_ ( .CLK(n22425), .D(n26684), .Q(n8180) );
  LATCH RN_reg_123_ ( .CLK(n22425), .D(n26719), .Q(n8179) );
  LATCH RN_reg_122_ ( .CLK(n22425), .D(n26768), .Q(n8178) );
  LATCH RN_reg_121_ ( .CLK(n22425), .D(n26825), .Q(n8177) );
  LATCH RN_reg_120_ ( .CLK(n22425), .D(n26883), .Q(n8176) );
  LATCH RN_reg_119_ ( .CLK(n22425), .D(n26952), .Q(n8175) );
  LATCH RN_reg_118_ ( .CLK(n22425), .D(n27030), .Q(n8174) );
  LATCH RN_reg_117_ ( .CLK(n22425), .D(n27125), .Q(n8173) );
  LATCH RN_reg_116_ ( .CLK(n22425), .D(n21336), .Q(n8172) );
  LATCH RN_reg_115_ ( .CLK(n22425), .D(n26579), .Q(n8171) );
  LATCH RN_reg_114_ ( .CLK(n22425), .D(n26601), .Q(n8170) );
  LATCH RN_reg_113_ ( .CLK(n22425), .D(n26627), .Q(n8169) );
  LATCH RN_reg_112_ ( .CLK(n22425), .D(n26653), .Q(n8168) );
  LATCH RN_reg_111_ ( .CLK(n22425), .D(n26685), .Q(n8167) );
  LATCH RN_reg_110_ ( .CLK(n22425), .D(n26720), .Q(n8166) );
  LATCH RN_reg_109_ ( .CLK(n22425), .D(n26769), .Q(n8165) );
  LATCH RN_reg_108_ ( .CLK(n22425), .D(n26826), .Q(n8164) );
  LATCH RN_reg_107_ ( .CLK(n22425), .D(n26884), .Q(n8163) );
  LATCH RN_reg_106_ ( .CLK(n22425), .D(n26953), .Q(n8162) );
  LATCH RN_reg_105_ ( .CLK(n22425), .D(n27031), .Q(n8161) );
  LATCH RN_reg_104_ ( .CLK(n22425), .D(n27126), .Q(n8160) );
  LATCH RN_reg_103_ ( .CLK(n22425), .D(n21333), .Q(n8159) );
  LATCH RN_reg_102_ ( .CLK(n22425), .D(n26582), .Q(n8158) );
  LATCH RN_reg_101_ ( .CLK(n22425), .D(n26604), .Q(n8157) );
  LATCH RN_reg_100_ ( .CLK(n22425), .D(n26630), .Q(n8156) );
  LATCH RN_reg_99_ ( .CLK(n22425), .D(n26656), .Q(n8155) );
  LATCH RN_reg_98_ ( .CLK(n22425), .D(n26688), .Q(n8154) );
  LATCH RN_reg_97_ ( .CLK(n22425), .D(n26723), .Q(n8153) );
  LATCH RN_reg_96_ ( .CLK(n22425), .D(n26772), .Q(n8152) );
  LATCH RN_reg_95_ ( .CLK(n22425), .D(n26829), .Q(n8151) );
  LATCH RN_reg_94_ ( .CLK(n22425), .D(n26887), .Q(n8150) );
  LATCH RN_reg_93_ ( .CLK(n22425), .D(n26956), .Q(n8149) );
  LATCH RN_reg_92_ ( .CLK(n22425), .D(n27034), .Q(n8148) );
  LATCH RN_reg_91_ ( .CLK(n22425), .D(n27129), .Q(n8147) );
  LATCH RN_reg_90_ ( .CLK(n22425), .D(n21330), .Q(n8146) );
  LATCH RN_reg_89_ ( .CLK(n22425), .D(n26583), .Q(n8145) );
  LATCH RN_reg_88_ ( .CLK(n22425), .D(n26605), .Q(n8144) );
  LATCH RN_reg_87_ ( .CLK(n22425), .D(n26631), .Q(n8143) );
  LATCH RN_reg_86_ ( .CLK(n22425), .D(n26657), .Q(n8142) );
  LATCH RN_reg_85_ ( .CLK(n22425), .D(n26689), .Q(n8141) );
  LATCH RN_reg_84_ ( .CLK(n22425), .D(n26724), .Q(n8140) );
  LATCH RN_reg_83_ ( .CLK(n22425), .D(n26773), .Q(n8139) );
  LATCH RN_reg_82_ ( .CLK(n22425), .D(n26830), .Q(n8138) );
  LATCH RN_reg_81_ ( .CLK(n22425), .D(n26888), .Q(n8137) );
  LATCH RN_reg_80_ ( .CLK(n22425), .D(n26957), .Q(n8136) );
  LATCH RN_reg_79_ ( .CLK(n22425), .D(n27035), .Q(n8135) );
  LATCH RN_reg_78_ ( .CLK(n22425), .D(n27130), .Q(n8134) );
  LATCH RN_reg_77_ ( .CLK(n22425), .D(n21327), .Q(n8133) );
  LATCH RN_reg_76_ ( .CLK(n22425), .D(n26584), .Q(n8132) );
  LATCH RN_reg_75_ ( .CLK(n22425), .D(n26606), .Q(n8131) );
  LATCH RN_reg_74_ ( .CLK(n22425), .D(n26632), .Q(n8130) );
  LATCH RN_reg_73_ ( .CLK(n22425), .D(n26658), .Q(n8129) );
  LATCH RN_reg_72_ ( .CLK(n22425), .D(n26690), .Q(n8128) );
  LATCH RN_reg_71_ ( .CLK(n22425), .D(n26725), .Q(n8127) );
  LATCH RN_reg_70_ ( .CLK(n22425), .D(n26774), .Q(n8126) );
  LATCH RN_reg_69_ ( .CLK(n22425), .D(n26831), .Q(n8125) );
  LATCH RN_reg_68_ ( .CLK(n22425), .D(n26889), .Q(n8124) );
  LATCH RN_reg_67_ ( .CLK(n22425), .D(n26958), .Q(n8123) );
  LATCH RN_reg_66_ ( .CLK(n22425), .D(n27036), .Q(n8122) );
  LATCH RN_reg_65_ ( .CLK(n22425), .D(n27131), .Q(n8121) );
  LATCH RN_reg_64_ ( .CLK(n22425), .D(n21326), .Q(n8120) );
  LATCH RN_reg_63_ ( .CLK(n22425), .D(n26585), .Q(n8119) );
  LATCH RN_reg_62_ ( .CLK(n22425), .D(n26607), .Q(n8118) );
  LATCH RN_reg_61_ ( .CLK(n22425), .D(n26633), .Q(n8117) );
  LATCH RN_reg_60_ ( .CLK(n22425), .D(n26659), .Q(n8116) );
  LATCH RN_reg_59_ ( .CLK(n22425), .D(n26691), .Q(n8115) );
  LATCH RN_reg_58_ ( .CLK(n22425), .D(n26726), .Q(n8114) );
  LATCH RN_reg_57_ ( .CLK(n22425), .D(n26775), .Q(n8113) );
  LATCH RN_reg_56_ ( .CLK(n22425), .D(n26832), .Q(n8112) );
  LATCH RN_reg_55_ ( .CLK(n22425), .D(n26890), .Q(n8111) );
  LATCH RN_reg_54_ ( .CLK(n22425), .D(n26959), .Q(n8110) );
  LATCH RN_reg_53_ ( .CLK(n22425), .D(n27037), .Q(n8109) );
  LATCH RN_reg_52_ ( .CLK(n22425), .D(n27132), .Q(n8108) );
  LATCH RN_reg_51_ ( .CLK(n22425), .D(n21321), .Q(n8107) );
  LATCH RN_reg_50_ ( .CLK(n22425), .D(n26586), .Q(n8106) );
  LATCH RN_reg_49_ ( .CLK(n22425), .D(n26608), .Q(n8105) );
  LATCH RN_reg_48_ ( .CLK(n22425), .D(n26634), .Q(n8104) );
  LATCH RN_reg_47_ ( .CLK(n22425), .D(n26660), .Q(n8103) );
  LATCH RN_reg_46_ ( .CLK(n22425), .D(n26692), .Q(n8102) );
  LATCH RN_reg_45_ ( .CLK(n22425), .D(n26727), .Q(n8101) );
  LATCH RN_reg_44_ ( .CLK(n22425), .D(n26776), .Q(n8100) );
  LATCH RN_reg_43_ ( .CLK(n22425), .D(n26833), .Q(n8099) );
  LATCH RN_reg_42_ ( .CLK(n22425), .D(n26891), .Q(n8098) );
  LATCH RN_reg_41_ ( .CLK(n22425), .D(n26960), .Q(n8097) );
  LATCH RN_reg_40_ ( .CLK(n22425), .D(n27038), .Q(n8096) );
  LATCH RN_reg_39_ ( .CLK(n22425), .D(n27133), .Q(n8095) );
  LATCH RN_reg_38_ ( .CLK(n22425), .D(n21320), .Q(n8094) );
  LATCH RN_reg_37_ ( .CLK(n22425), .D(n26587), .Q(n8093) );
  LATCH RN_reg_36_ ( .CLK(n22425), .D(n26609), .Q(n8092) );
  LATCH RN_reg_35_ ( .CLK(n22425), .D(n26635), .Q(n8091) );
  LATCH RN_reg_34_ ( .CLK(n22425), .D(n26661), .Q(n8090) );
  LATCH RN_reg_33_ ( .CLK(n22425), .D(n26693), .Q(n8089) );
  LATCH RN_reg_32_ ( .CLK(n22425), .D(n26728), .Q(n8088) );
  LATCH RN_reg_31_ ( .CLK(n22425), .D(n26777), .Q(n8087) );
  LATCH RN_reg_30_ ( .CLK(n22425), .D(n26834), .Q(n8086) );
  LATCH RN_reg_29_ ( .CLK(n22425), .D(n26892), .Q(n8085) );
  LATCH RN_reg_28_ ( .CLK(n22425), .D(n26961), .Q(n8084) );
  LATCH RN_reg_27_ ( .CLK(n22425), .D(n27039), .Q(n8083) );
  LATCH RN_reg_26_ ( .CLK(n22425), .D(n27134), .Q(n8082) );
  LATCH RN_reg_25_ ( .CLK(n22425), .D(n26611), .Q(n8081) );
  LATCH RN_reg_24_ ( .CLK(n22425), .D(n26637), .Q(n8080) );
  LATCH RN_reg_23_ ( .CLK(n22425), .D(n26663), .Q(n8079) );
  LATCH RN_reg_22_ ( .CLK(n22425), .D(n26695), .Q(n8078) );
  LATCH RN_reg_21_ ( .CLK(n22425), .D(n26730), .Q(n8077) );
  LATCH RN_reg_20_ ( .CLK(n22425), .D(n26778), .Q(n8076) );
  LATCH RN_reg_19_ ( .CLK(n22425), .D(n26835), .Q(n8075) );
  LATCH RN_reg_18_ ( .CLK(n22425), .D(n26893), .Q(n8074) );
  LATCH RN_reg_17_ ( .CLK(n22425), .D(n27135), .Q(n8073) );
  LATCH RN_reg_16_ ( .CLK(n22425), .D(n27136), .Q(n8072) );
  LATCH RN_reg_15_ ( .CLK(n22425), .D(n27137), .Q(n8071) );
  LATCH RN_reg_14_ ( .CLK(n22425), .D(n26962), .Q(n8070) );
  LATCH RN_reg_13_ ( .CLK(n22425), .D(n27040), .Q(n8069) );
  LATCH RN_reg_12_ ( .CLK(n22425), .D(n26779), .Q(n8068) );
  LATCH RN_reg_11_ ( .CLK(n22425), .D(n26836), .Q(n8067) );
  LATCH RN_reg_10_ ( .CLK(n22425), .D(n26894), .Q(n8066) );
  LATCH RN_reg_9_ ( .CLK(n22425), .D(n26963), .Q(n8065) );
  LATCH RN_reg_8_ ( .CLK(n22425), .D(n27138), .Q(n8064) );
  LATCH RN_reg_7_ ( .CLK(n22425), .D(n27139), .Q(n8063) );
  LATCH RN_reg_6_ ( .CLK(n22425), .D(n27041), .Q(n8062) );
  LATCH RN_reg_5_ ( .CLK(n22425), .D(n26729), .Q(n8061) );
  LATCH RN_reg_4_ ( .CLK(n22425), .D(n21319), .Q(n8060) );
  LATCH RN_reg_3_ ( .CLK(n22425), .D(n26636), .Q(n8059) );
  LATCH RN_reg_2_ ( .CLK(n22425), .D(n26694), .Q(n8058) );
  LATCH RN_reg_1_ ( .CLK(n22425), .D(n26662), .Q(n8057) );
  LATCH RN_reg_0_ ( .CLK(n22425), .D(n26610), .Q(n8056) );
  LATCH we_reg ( .CLK(n22324), .D(net96340), .Q(we) );
  LATCH loc_s2_reg_0_ ( .CLK(n22637), .D(n13703), .Q(loc_s2[0]) );
  LATCH loc_s2_reg_1_ ( .CLK(n22637), .D(n13704), .Q(loc_s2[1]) );
  LATCH loc_s2_reg_2_ ( .CLK(n22637), .D(n13705), .Q(loc_s2[2]) );
  LATCH loc_s2_reg_3_ ( .CLK(n22637), .D(n13706), .Q(loc_s2[3]) );
  LATCH loc_s2_reg_4_ ( .CLK(n22637), .D(n23085), .Q(loc_s2[4]) );
  LATCH loc_s2_reg_5_ ( .CLK(n22637), .D(n24982), .Q(loc_s2[5]) );
  LATCH invdirect_s2_reg_0_ ( .CLK(n22637), .D(n27181), .Q(invdirect_s2[0]) );
  LATCH invdirect_s2_reg_1_ ( .CLK(n22637), .D(n24927), .Q(invdirect_s2[1]) );
  LATCH invdirect_s2_reg_2_ ( .CLK(n22637), .D(n34503), .Q(invdirect_s2[2]) );
  LATCH oc_reg_0_ ( .CLK(n22426), .D(n21312), .Q(oc[0]) );
  LATCH oc_reg_29_ ( .CLK(n22426), .D(n21311), .Q(oc[29]) );
  LATCH oc_reg_1_ ( .CLK(n22426), .D(n23628), .Q(oc[1]) );
  LATCH oc_reg_2_ ( .CLK(n22426), .D(n21310), .Q(oc[2]) );
  LATCH oc_reg_3_ ( .CLK(n22426), .D(n21309), .Q(oc[3]) );
  LATCH oc_reg_4_ ( .CLK(n22426), .D(n26780), .Q(oc[4]) );
  LATCH oc_reg_5_ ( .CLK(n22426), .D(n21308), .Q(oc[5]) );
  LATCH oc_reg_6_ ( .CLK(n22426), .D(n23627), .Q(oc[6]) );
  LATCH oc_reg_7_ ( .CLK(n22426), .D(n23626), .Q(oc[7]) );
  LATCH oc_reg_8_ ( .CLK(n22426), .D(n21307), .Q(oc[8]) );
  LATCH oc_reg_9_ ( .CLK(n22426), .D(n21306), .Q(oc[9]) );
  LATCH oc_reg_10_ ( .CLK(n22426), .D(n21305), .Q(oc[10]) );
  LATCH oc_reg_11_ ( .CLK(n22426), .D(n21304), .Q(oc[11]) );
  LATCH oc_reg_12_ ( .CLK(n22426), .D(n21303), .Q(oc[12]) );
  LATCH oc_reg_13_ ( .CLK(n22426), .D(n21302), .Q(oc[13]) );
  LATCH oc_reg_14_ ( .CLK(n22426), .D(n21301), .Q(oc[14]) );
  LATCH oc_reg_15_ ( .CLK(n22426), .D(n21300), .Q(oc[15]) );
  LATCH oc_reg_16_ ( .CLK(n22426), .D(n21299), .Q(oc[16]) );
  LATCH oc_reg_17_ ( .CLK(n22426), .D(n21298), .Q(oc[17]) );
  LATCH oc_reg_18_ ( .CLK(n22426), .D(net146640), .Q(oc[18]) );
  LATCH oc_reg_19_ ( .CLK(n22426), .D(n21297), .Q(oc[19]) );
  LATCH oc_reg_20_ ( .CLK(n22426), .D(n21296), .Q(oc[20]) );
  LATCH oc_reg_21_ ( .CLK(n22426), .D(n21295), .Q(oc[21]) );
  LATCH oc_reg_22_ ( .CLK(n22426), .D(n21294), .Q(oc[22]) );
  LATCH oc_reg_23_ ( .CLK(n22426), .D(n21293), .Q(oc[23]) );
  LATCH oc_reg_24_ ( .CLK(n22426), .D(n21292), .Q(oc[24]) );
  LATCH oc_reg_25_ ( .CLK(n22426), .D(n21291), .Q(oc[25]) );
  LATCH oc_reg_26_ ( .CLK(n22426), .D(n21290), .Q(oc[26]) );
  LATCH oc_reg_27_ ( .CLK(n22426), .D(n21289), .Q(oc[27]) );
  LATCH oc_reg_28_ ( .CLK(n22426), .D(n21288), .Q(oc[28]) );
  LATCH Setup_reg_0_ ( .CLK(n22328), .D(n27122), .Q(Setup[0]) );
  LATCH Setup_reg_1_ ( .CLK(n22328), .D(n26949), .Q(Setup[1]) );
  LATCH S_reg_0_ ( .CLK(n22626), .D(data_in[0]), .Q(S[0]) );
  LATCH S_reg_1_ ( .CLK(n22626), .D(data_in[1]), .Q(S[1]) );
  LATCH S_reg_2_ ( .CLK(n22626), .D(data_in[2]), .Q(S[2]) );
  LATCH S_reg_3_ ( .CLK(n22626), .D(data_in[3]), .Q(S[3]) );
  LATCH S_reg_4_ ( .CLK(n22626), .D(data_in[4]), .Q(S[4]) );
  LATCH S_reg_5_ ( .CLK(n22626), .D(data_in[5]), .Q(S[5]) );
  LATCH wS_reg ( .CLK(n22428), .D(net96340), .Q(wS) );
  LATCH D_reg ( .CLK(n22326), .D(net96340), .Q(D) );
  LATCH wT_reg ( .CLK(n22427), .D(net96340), .Q(wT) );
  LATCH location_reg_0_ ( .CLK(n22632), .D(n20534), .Q(n2251) );
  LATCH location_reg_1_ ( .CLK(n22632), .D(n21287), .Q(n2252) );
  LATCH cs_reg ( .CLK(n22323), .D(net96340), .Q(cs) );
  LATCH T_reg_1_ ( .CLK(n22627), .D(data_in[1]), .Q(T[1]) );
  LATCH T_reg_2_ ( .CLK(n22627), .D(data_in[2]), .Q(T[2]) );
  LATCH T_reg_3_ ( .CLK(n22627), .D(data_in[3]), .Q(T[3]) );
  LATCH T_reg_4_ ( .CLK(n22627), .D(data_in[4]), .Q(T[4]) );
  LATCH T_reg_5_ ( .CLK(n22627), .D(data_in[5]), .Q(T[5]) );
  LATCH RO_reg_126_ ( .CLK(n22393), .D(n21518), .Q(n3228) );
  LATCH RO_reg_2_ ( .CLK(n22330), .D(n21331), .Q(n3104) );
  LATCH RO_reg_3_ ( .CLK(n22330), .D(n21332), .Q(n3105) );
  LATCH RO_reg_4_ ( .CLK(n22331), .D(n21334), .Q(n3106) );
  LATCH RO_reg_5_ ( .CLK(n22331), .D(n21335), .Q(n3107) );
  LATCH RO_reg_6_ ( .CLK(n22332), .D(n21337), .Q(n3108) );
  LATCH RO_reg_7_ ( .CLK(n22332), .D(n21338), .Q(n3109) );
  LATCH RO_reg_8_ ( .CLK(n22333), .D(n21286), .Q(n3110) );
  LATCH RO_reg_9_ ( .CLK(n22333), .D(n21285), .Q(n3111) );
  LATCH RO_reg_10_ ( .CLK(n22334), .D(n21343), .Q(n3112) );
  LATCH RO_reg_11_ ( .CLK(n22334), .D(n21344), .Q(n3113) );
  LATCH RO_reg_12_ ( .CLK(n22335), .D(n21346), .Q(n3114) );
  LATCH RO_reg_13_ ( .CLK(n22335), .D(n21347), .Q(n3115) );
  LATCH RO_reg_14_ ( .CLK(n22336), .D(n21284), .Q(n3116) );
  LATCH RO_reg_15_ ( .CLK(n22336), .D(n21283), .Q(n3117) );
  LATCH RO_reg_16_ ( .CLK(n22337), .D(n21352), .Q(n3118) );
  LATCH RO_reg_17_ ( .CLK(n22337), .D(n21353), .Q(n3119) );
  LATCH RO_reg_18_ ( .CLK(n22338), .D(n21355), .Q(n3120) );
  LATCH RO_reg_19_ ( .CLK(n22338), .D(n21356), .Q(n3121) );
  LATCH RO_reg_20_ ( .CLK(n22339), .D(n21282), .Q(n3122) );
  LATCH RO_reg_21_ ( .CLK(n22339), .D(n21281), .Q(n3123) );
  LATCH RO_reg_22_ ( .CLK(n22340), .D(n21361), .Q(n3124) );
  LATCH RO_reg_23_ ( .CLK(n22340), .D(n21362), .Q(n3125) );
  LATCH RO_reg_24_ ( .CLK(n22341), .D(n21364), .Q(n3126) );
  LATCH RO_reg_25_ ( .CLK(n22341), .D(n21365), .Q(n3127) );
  LATCH RO_reg_26_ ( .CLK(n22342), .D(n21280), .Q(n3128) );
  LATCH RO_reg_27_ ( .CLK(n22342), .D(n21279), .Q(n3129) );
  LATCH RO_reg_28_ ( .CLK(n22343), .D(n21370), .Q(n3130) );
  LATCH RO_reg_29_ ( .CLK(n22343), .D(n21371), .Q(n3131) );
  LATCH RO_reg_30_ ( .CLK(n22344), .D(n21373), .Q(n3132) );
  LATCH RO_reg_31_ ( .CLK(n22344), .D(n21374), .Q(n3133) );
  LATCH RO_reg_32_ ( .CLK(n22345), .D(n21278), .Q(n3134) );
  LATCH RO_reg_33_ ( .CLK(n22345), .D(n21277), .Q(n3135) );
  LATCH RO_reg_34_ ( .CLK(n22346), .D(n21379), .Q(n3136) );
  LATCH RO_reg_35_ ( .CLK(n22346), .D(n21380), .Q(n3137) );
  LATCH RO_reg_36_ ( .CLK(n22347), .D(n21382), .Q(n3138) );
  LATCH RO_reg_37_ ( .CLK(n22347), .D(n21383), .Q(n3139) );
  LATCH RO_reg_38_ ( .CLK(n22348), .D(n21276), .Q(n3140) );
  LATCH RO_reg_39_ ( .CLK(n22348), .D(n21275), .Q(n3141) );
  LATCH RO_reg_40_ ( .CLK(n22349), .D(n21388), .Q(n3142) );
  LATCH RO_reg_41_ ( .CLK(n22349), .D(n21389), .Q(n3143) );
  LATCH RO_reg_42_ ( .CLK(n22350), .D(n21391), .Q(n3144) );
  LATCH RO_reg_43_ ( .CLK(n22350), .D(n21392), .Q(n3145) );
  LATCH RO_reg_44_ ( .CLK(n22351), .D(n21274), .Q(n3146) );
  LATCH RO_reg_45_ ( .CLK(n22351), .D(n21273), .Q(n3147) );
  LATCH RO_reg_46_ ( .CLK(n22352), .D(n21397), .Q(n3148) );
  LATCH RO_reg_47_ ( .CLK(n22352), .D(n21398), .Q(n3149) );
  LATCH RO_reg_48_ ( .CLK(n22353), .D(n21400), .Q(n3150) );
  LATCH RO_reg_49_ ( .CLK(n22353), .D(n21401), .Q(n3151) );
  LATCH RO_reg_50_ ( .CLK(n22354), .D(n21272), .Q(n3152) );
  LATCH RO_reg_51_ ( .CLK(n22354), .D(n21271), .Q(n3153) );
  LATCH RO_reg_52_ ( .CLK(n22355), .D(n21406), .Q(n3154) );
  LATCH RO_reg_53_ ( .CLK(n22355), .D(n21407), .Q(n3155) );
  LATCH RO_reg_54_ ( .CLK(n22356), .D(n21409), .Q(n3156) );
  LATCH RO_reg_55_ ( .CLK(n22356), .D(n21410), .Q(n3157) );
  LATCH RO_reg_56_ ( .CLK(n22357), .D(n21270), .Q(n3158) );
  LATCH RO_reg_57_ ( .CLK(n22357), .D(n21269), .Q(n3159) );
  LATCH RO_reg_58_ ( .CLK(n22358), .D(n21415), .Q(n3160) );
  LATCH RO_reg_59_ ( .CLK(n22358), .D(n21416), .Q(n3161) );
  LATCH RO_reg_60_ ( .CLK(n22359), .D(n21418), .Q(n3162) );
  LATCH RO_reg_61_ ( .CLK(n22359), .D(n21419), .Q(n3163) );
  LATCH RO_reg_62_ ( .CLK(n22360), .D(n21268), .Q(n3164) );
  LATCH RO_reg_63_ ( .CLK(n22360), .D(n21267), .Q(n3165) );
  LATCH RO_reg_64_ ( .CLK(n22361), .D(n21424), .Q(n3166) );
  LATCH RO_reg_65_ ( .CLK(n22361), .D(n21425), .Q(n3167) );
  LATCH RO_reg_66_ ( .CLK(n22362), .D(n21427), .Q(n3168) );
  LATCH RO_reg_67_ ( .CLK(n22362), .D(n21428), .Q(n3169) );
  LATCH RO_reg_68_ ( .CLK(n22363), .D(n21266), .Q(n3170) );
  LATCH RO_reg_69_ ( .CLK(n22363), .D(n21265), .Q(n3171) );
  LATCH RO_reg_70_ ( .CLK(n22364), .D(n21433), .Q(n3172) );
  LATCH RO_reg_71_ ( .CLK(n22364), .D(n21434), .Q(n3173) );
  LATCH RO_reg_72_ ( .CLK(n22365), .D(n21436), .Q(n3174) );
  LATCH RO_reg_73_ ( .CLK(n22365), .D(n21437), .Q(n3175) );
  LATCH RO_reg_74_ ( .CLK(n22366), .D(n21264), .Q(n3176) );
  LATCH RO_reg_75_ ( .CLK(n22366), .D(n21263), .Q(n3177) );
  LATCH RO_reg_76_ ( .CLK(n22367), .D(n21442), .Q(n3178) );
  LATCH RO_reg_77_ ( .CLK(n22367), .D(n21443), .Q(n3179) );
  LATCH RO_reg_78_ ( .CLK(n22368), .D(n21445), .Q(n3180) );
  LATCH RO_reg_79_ ( .CLK(n22368), .D(n21446), .Q(n3181) );
  LATCH RO_reg_80_ ( .CLK(n22369), .D(n21262), .Q(n3182) );
  LATCH RO_reg_81_ ( .CLK(n22369), .D(n21261), .Q(n3183) );
  LATCH RO_reg_82_ ( .CLK(n22370), .D(n21451), .Q(n3184) );
  LATCH RO_reg_83_ ( .CLK(n22370), .D(n21452), .Q(n3185) );
  LATCH RO_reg_84_ ( .CLK(n22371), .D(n21454), .Q(n3186) );
  LATCH RO_reg_85_ ( .CLK(n22371), .D(n21455), .Q(n3187) );
  LATCH RO_reg_86_ ( .CLK(n22372), .D(n21260), .Q(n3188) );
  LATCH RO_reg_87_ ( .CLK(n22372), .D(n21259), .Q(n3189) );
  LATCH RO_reg_88_ ( .CLK(n22373), .D(n21460), .Q(n3190) );
  LATCH RO_reg_89_ ( .CLK(n22373), .D(n21461), .Q(n3191) );
  LATCH RO_reg_90_ ( .CLK(n22374), .D(n21463), .Q(n3192) );
  LATCH RO_reg_91_ ( .CLK(n22374), .D(n21464), .Q(n3193) );
  LATCH RO_reg_92_ ( .CLK(n22376), .D(n21258), .Q(n3194) );
  LATCH RO_reg_93_ ( .CLK(n22376), .D(n21257), .Q(n3195) );
  LATCH RO_reg_94_ ( .CLK(n22377), .D(n21470), .Q(n3196) );
  LATCH RO_reg_95_ ( .CLK(n22377), .D(n21471), .Q(n3197) );
  LATCH RO_reg_96_ ( .CLK(n22378), .D(n21473), .Q(n3198) );
  LATCH RO_reg_97_ ( .CLK(n22378), .D(n21474), .Q(n3199) );
  LATCH RO_reg_98_ ( .CLK(n22379), .D(n21476), .Q(n3200) );
  LATCH RO_reg_99_ ( .CLK(n22379), .D(n21477), .Q(n3201) );
  LATCH RO_reg_100_ ( .CLK(n22380), .D(n21479), .Q(n3202) );
  LATCH RO_reg_101_ ( .CLK(n22380), .D(n21480), .Q(n3203) );
  LATCH RO_reg_102_ ( .CLK(n22381), .D(n21482), .Q(n3204) );
  LATCH RO_reg_103_ ( .CLK(n22381), .D(n21483), .Q(n3205) );
  LATCH RO_reg_104_ ( .CLK(n22382), .D(n21256), .Q(n3206) );
  LATCH RO_reg_105_ ( .CLK(n22382), .D(n21255), .Q(n3207) );
  LATCH RO_reg_106_ ( .CLK(n22383), .D(n21488), .Q(n3208) );
  LATCH RO_reg_107_ ( .CLK(n22383), .D(n21489), .Q(n3209) );
  LATCH RO_reg_108_ ( .CLK(n22384), .D(n21491), .Q(n3210) );
  LATCH RO_reg_109_ ( .CLK(n22384), .D(n21492), .Q(n3211) );
  LATCH RO_reg_110_ ( .CLK(n22385), .D(n21254), .Q(n3212) );
  LATCH RO_reg_111_ ( .CLK(n22385), .D(n21253), .Q(n3213) );
  LATCH RO_reg_112_ ( .CLK(n22386), .D(n21497), .Q(n3214) );
  LATCH RO_reg_113_ ( .CLK(n22386), .D(n21498), .Q(n3215) );
  LATCH RO_reg_114_ ( .CLK(n22387), .D(n21500), .Q(n3216) );
  LATCH RO_reg_115_ ( .CLK(n22387), .D(n21501), .Q(n3217) );
  LATCH RO_reg_116_ ( .CLK(n22388), .D(n21252), .Q(n3218) );
  LATCH RO_reg_117_ ( .CLK(n22388), .D(n21251), .Q(n3219) );
  LATCH RO_reg_118_ ( .CLK(n22389), .D(n21506), .Q(n3220) );
  LATCH RO_reg_119_ ( .CLK(n22389), .D(n21507), .Q(n3221) );
  LATCH RO_reg_120_ ( .CLK(n22390), .D(n21509), .Q(n3222) );
  LATCH RO_reg_121_ ( .CLK(n22390), .D(n21510), .Q(n3223) );
  LATCH RO_reg_122_ ( .CLK(n22391), .D(n21250), .Q(n3224) );
  LATCH RO_reg_123_ ( .CLK(n22391), .D(n21249), .Q(n3225) );
  LATCH RO_reg_124_ ( .CLK(n22392), .D(n21515), .Q(n3226) );
  LATCH RO_reg_125_ ( .CLK(n22392), .D(n21516), .Q(n3227) );
  LATCH RO_reg_127_ ( .CLK(n22393), .D(n21519), .Q(n3229) );
  LATCH RO_reg_128_ ( .CLK(n22394), .D(n21248), .Q(n3230) );
  LATCH RO_reg_129_ ( .CLK(n22394), .D(n34459), .Q(n3231) );
  LATCH RO_reg_130_ ( .CLK(n22395), .D(n34492), .Q(n3232) );
  LATCH RO_reg_131_ ( .CLK(n22395), .D(n34491), .Q(n3233) );
  LATCH RO_reg_132_ ( .CLK(n22396), .D(n34490), .Q(n3234) );
  LATCH RO_reg_133_ ( .CLK(n22396), .D(n34489), .Q(n3235) );
  LATCH RO_reg_134_ ( .CLK(n22397), .D(n34458), .Q(n3236) );
  LATCH RO_reg_135_ ( .CLK(n22397), .D(n34457), .Q(n3237) );
  LATCH RO_reg_136_ ( .CLK(n22398), .D(n34488), .Q(n3238) );
  LATCH RO_reg_137_ ( .CLK(n22398), .D(n34487), .Q(n3239) );
  LATCH RO_reg_138_ ( .CLK(n22399), .D(n34486), .Q(n3240) );
  LATCH RO_reg_139_ ( .CLK(n22399), .D(n34485), .Q(n3241) );
  LATCH RO_reg_140_ ( .CLK(n22400), .D(n34456), .Q(n3242) );
  LATCH RO_reg_141_ ( .CLK(n22400), .D(n34455), .Q(n3243) );
  LATCH RO_reg_142_ ( .CLK(n22401), .D(n34484), .Q(n3244) );
  LATCH RO_reg_143_ ( .CLK(n22401), .D(n34483), .Q(n3245) );
  LATCH RO_reg_144_ ( .CLK(n22402), .D(n34482), .Q(n3246) );
  LATCH RO_reg_145_ ( .CLK(n22402), .D(n34481), .Q(n3247) );
  LATCH RO_reg_146_ ( .CLK(n22403), .D(n34454), .Q(n3248) );
  LATCH RO_reg_147_ ( .CLK(n22403), .D(n34453), .Q(n3249) );
  LATCH RO_reg_148_ ( .CLK(n22404), .D(n34480), .Q(n3250) );
  LATCH RO_reg_149_ ( .CLK(n22404), .D(n34479), .Q(n3251) );
  LATCH RO_reg_150_ ( .CLK(n22405), .D(n34478), .Q(n3252) );
  LATCH RO_reg_151_ ( .CLK(n22405), .D(n34477), .Q(n3253) );
  LATCH RO_reg_152_ ( .CLK(n22406), .D(n34452), .Q(n3254) );
  LATCH RO_reg_153_ ( .CLK(n22406), .D(n34451), .Q(n3255) );
  LATCH RO_reg_154_ ( .CLK(n22407), .D(n34476), .Q(n3256) );
  LATCH RO_reg_155_ ( .CLK(n22407), .D(n34475), .Q(n3257) );
  LATCH RO_reg_156_ ( .CLK(n22408), .D(n34474), .Q(n3258) );
  LATCH RO_reg_157_ ( .CLK(n22408), .D(n34473), .Q(n3259) );
  LATCH RO_reg_158_ ( .CLK(n22409), .D(n34450), .Q(n3260) );
  LATCH RO_reg_159_ ( .CLK(n22409), .D(n34449), .Q(n3261) );
  LATCH RO_reg_160_ ( .CLK(n22410), .D(n34472), .Q(n3262) );
  LATCH RO_reg_161_ ( .CLK(n22410), .D(n34471), .Q(n3263) );
  LATCH RO_reg_162_ ( .CLK(n22411), .D(n34470), .Q(n3264) );
  LATCH RO_reg_163_ ( .CLK(n22411), .D(n34469), .Q(n3265) );
  LATCH RO_reg_164_ ( .CLK(n22412), .D(n34448), .Q(n3266) );
  LATCH RO_reg_165_ ( .CLK(n22412), .D(n34447), .Q(n3267) );
  LATCH RO_reg_166_ ( .CLK(n22413), .D(n34468), .Q(n3268) );
  LATCH RO_reg_167_ ( .CLK(n22413), .D(n34467), .Q(n3269) );
  LATCH RO_reg_168_ ( .CLK(n22414), .D(n34466), .Q(n3270) );
  LATCH RO_reg_169_ ( .CLK(n22414), .D(n34465), .Q(n3271) );
  LATCH RO_reg_170_ ( .CLK(n22415), .D(n34446), .Q(n3272) );
  LATCH RO_reg_171_ ( .CLK(n22415), .D(n34445), .Q(n3273) );
  LATCH RO_reg_172_ ( .CLK(n22416), .D(n34464), .Q(n3274) );
  LATCH RO_reg_173_ ( .CLK(n22416), .D(n34463), .Q(n3275) );
  LATCH RO_reg_174_ ( .CLK(n22417), .D(n34462), .Q(RO[174]) );
  LATCH RO_reg_175_ ( .CLK(n22417), .D(n34461), .Q(RO[175]) );
  LATCH RO_reg_176_ ( .CLK(n22418), .D(n34444), .Q(RO[176]) );
  LATCH locTrig_reg_1_ ( .CLK(n22431), .D(n21176), .Q(locTrig[1]) );
  LATCH direction_lee_reg_1_ ( .CLK(n22636), .D(n24981), .Q(direction_lee[1])
         );
  LATCH locTrig_reg_3_ ( .CLK(n22433), .D(n21247), .Q(locTrig[3]) );
  LATCH direction_lee_reg_0_ ( .CLK(n22636), .D(n22881), .Q(direction_lee[0])
         );
  LATCH pLoc_reg_1_ ( .CLK(n22629), .D(n11045), .Q(pLoc[1]) );
  LATCH grid_reg_63__4_ ( .CLK(n22625), .D(n29458), .Q(grid[382]) );
  LATCH grid_reg_63__5_ ( .CLK(n22625), .D(n29449), .Q(grid[383]) );
  LATCH grid_reg_62__4_ ( .CLK(n22622), .D(n29458), .Q(grid[376]) );
  LATCH grid_reg_62__5_ ( .CLK(n22622), .D(n29449), .Q(grid[377]) );
  LATCH grid_reg_61__4_ ( .CLK(n22619), .D(n29458), .Q(grid[370]) );
  LATCH grid_reg_61__5_ ( .CLK(n22619), .D(n29449), .Q(grid[371]) );
  LATCH grid_reg_60__4_ ( .CLK(n22616), .D(n29458), .Q(grid[364]) );
  LATCH grid_reg_60__5_ ( .CLK(n22616), .D(n29449), .Q(grid[365]) );
  LATCH grid_reg_59__4_ ( .CLK(n22613), .D(n29457), .Q(grid[358]) );
  LATCH grid_reg_59__5_ ( .CLK(n22613), .D(n29448), .Q(grid[359]) );
  LATCH grid_reg_58__4_ ( .CLK(n22610), .D(n29457), .Q(grid[352]) );
  LATCH grid_reg_58__5_ ( .CLK(n22610), .D(n29448), .Q(grid[353]) );
  LATCH grid_reg_57__4_ ( .CLK(n22607), .D(n29457), .Q(grid[346]) );
  LATCH grid_reg_57__5_ ( .CLK(n22607), .D(n29448), .Q(grid[347]) );
  LATCH grid_reg_56__4_ ( .CLK(n22604), .D(n29457), .Q(grid[340]) );
  LATCH grid_reg_56__5_ ( .CLK(n22604), .D(n29448), .Q(grid[341]) );
  LATCH grid_reg_55__4_ ( .CLK(n22601), .D(n29457), .Q(grid[334]) );
  LATCH grid_reg_55__5_ ( .CLK(n22601), .D(n29448), .Q(grid[335]) );
  LATCH grid_reg_54__4_ ( .CLK(n22598), .D(n29457), .Q(grid[328]) );
  LATCH grid_reg_54__5_ ( .CLK(n22598), .D(n29448), .Q(grid[329]) );
  LATCH grid_reg_53__4_ ( .CLK(n22595), .D(n29457), .Q(grid[322]) );
  LATCH grid_reg_53__5_ ( .CLK(n22595), .D(n29448), .Q(grid[323]) );
  LATCH grid_reg_52__4_ ( .CLK(n22592), .D(n29457), .Q(grid[316]) );
  LATCH grid_reg_52__5_ ( .CLK(n22592), .D(n29448), .Q(grid[317]) );
  LATCH grid_reg_51__4_ ( .CLK(n22589), .D(n29457), .Q(grid[310]) );
  LATCH grid_reg_51__5_ ( .CLK(n22589), .D(n29448), .Q(grid[311]) );
  LATCH grid_reg_50__4_ ( .CLK(n22586), .D(n29457), .Q(grid[304]) );
  LATCH grid_reg_50__5_ ( .CLK(n22586), .D(n29448), .Q(grid[305]) );
  LATCH grid_reg_49__4_ ( .CLK(n22583), .D(n29457), .Q(grid[298]) );
  LATCH grid_reg_49__5_ ( .CLK(n22583), .D(n29448), .Q(grid[299]) );
  LATCH grid_reg_48__4_ ( .CLK(n22580), .D(n29457), .Q(grid[292]) );
  LATCH grid_reg_48__5_ ( .CLK(n22580), .D(n29448), .Q(grid[293]) );
  LATCH grid_reg_47__4_ ( .CLK(n22577), .D(n29456), .Q(grid[286]) );
  LATCH grid_reg_47__5_ ( .CLK(n22577), .D(n29447), .Q(grid[287]) );
  LATCH grid_reg_46__4_ ( .CLK(n22574), .D(n29456), .Q(grid[280]) );
  LATCH grid_reg_46__5_ ( .CLK(n22574), .D(n29447), .Q(grid[281]) );
  LATCH grid_reg_45__4_ ( .CLK(n22571), .D(n29456), .Q(grid[274]) );
  LATCH grid_reg_45__5_ ( .CLK(n22571), .D(n29447), .Q(grid[275]) );
  LATCH grid_reg_44__4_ ( .CLK(n22568), .D(n29456), .Q(grid[268]) );
  LATCH grid_reg_44__5_ ( .CLK(n22568), .D(n29447), .Q(grid[269]) );
  LATCH grid_reg_43__4_ ( .CLK(n22565), .D(n29456), .Q(grid[262]) );
  LATCH grid_reg_43__5_ ( .CLK(n22565), .D(n29447), .Q(grid[263]) );
  LATCH grid_reg_42__4_ ( .CLK(n22562), .D(n29456), .Q(grid[256]) );
  LATCH grid_reg_42__5_ ( .CLK(n22562), .D(n29447), .Q(grid[257]) );
  LATCH grid_reg_41__4_ ( .CLK(n22559), .D(n29456), .Q(grid[250]) );
  LATCH grid_reg_41__5_ ( .CLK(n22559), .D(n29447), .Q(grid[251]) );
  LATCH grid_reg_40__4_ ( .CLK(n22556), .D(n29456), .Q(grid[244]) );
  LATCH grid_reg_40__5_ ( .CLK(n22556), .D(n29447), .Q(grid[245]) );
  LATCH grid_reg_39__4_ ( .CLK(n22553), .D(n29456), .Q(grid[238]) );
  LATCH grid_reg_39__5_ ( .CLK(n22553), .D(n29447), .Q(grid[239]) );
  LATCH grid_reg_38__4_ ( .CLK(n22550), .D(n29456), .Q(grid[232]) );
  LATCH grid_reg_38__5_ ( .CLK(n22550), .D(n29447), .Q(grid[233]) );
  LATCH grid_reg_37__4_ ( .CLK(n22547), .D(n29456), .Q(grid[226]) );
  LATCH grid_reg_37__5_ ( .CLK(n22547), .D(n29447), .Q(grid[227]) );
  LATCH grid_reg_36__4_ ( .CLK(n22544), .D(n29456), .Q(grid[220]) );
  LATCH grid_reg_36__5_ ( .CLK(n22544), .D(n29447), .Q(grid[221]) );
  LATCH grid_reg_35__4_ ( .CLK(n22541), .D(n29455), .Q(grid[214]) );
  LATCH grid_reg_35__5_ ( .CLK(n22541), .D(n29446), .Q(grid[215]) );
  LATCH grid_reg_34__4_ ( .CLK(n22538), .D(n29455), .Q(grid[208]) );
  LATCH grid_reg_34__5_ ( .CLK(n22538), .D(n29446), .Q(grid[209]) );
  LATCH grid_reg_33__4_ ( .CLK(n22535), .D(n29455), .Q(grid[202]) );
  LATCH grid_reg_33__5_ ( .CLK(n22535), .D(n29446), .Q(grid[203]) );
  LATCH grid_reg_32__4_ ( .CLK(n22532), .D(n29455), .Q(grid[196]) );
  LATCH grid_reg_32__5_ ( .CLK(n22532), .D(n29446), .Q(grid[197]) );
  LATCH grid_reg_31__4_ ( .CLK(n22529), .D(n29455), .Q(grid[190]) );
  LATCH grid_reg_31__5_ ( .CLK(n22529), .D(n29446), .Q(grid[191]) );
  LATCH grid_reg_30__4_ ( .CLK(n22526), .D(n29455), .Q(grid[184]) );
  LATCH grid_reg_30__5_ ( .CLK(n22526), .D(n29446), .Q(grid[185]) );
  LATCH grid_reg_29__4_ ( .CLK(n22523), .D(n29455), .Q(grid[178]) );
  LATCH grid_reg_29__5_ ( .CLK(n22523), .D(n29446), .Q(grid[179]) );
  LATCH grid_reg_28__4_ ( .CLK(n22520), .D(n29455), .Q(grid[172]) );
  LATCH grid_reg_28__5_ ( .CLK(n22520), .D(n29446), .Q(grid[173]) );
  LATCH grid_reg_27__4_ ( .CLK(n22517), .D(n29455), .Q(grid[166]) );
  LATCH grid_reg_27__5_ ( .CLK(n22517), .D(n29446), .Q(grid[167]) );
  LATCH grid_reg_26__4_ ( .CLK(n22514), .D(n29455), .Q(grid[160]) );
  LATCH grid_reg_26__5_ ( .CLK(n22514), .D(n29446), .Q(grid[161]) );
  LATCH grid_reg_25__4_ ( .CLK(n22511), .D(n29455), .Q(grid[154]) );
  LATCH grid_reg_25__5_ ( .CLK(n22511), .D(n29446), .Q(grid[155]) );
  LATCH grid_reg_24__4_ ( .CLK(n22508), .D(n29455), .Q(grid[148]) );
  LATCH grid_reg_24__5_ ( .CLK(n22508), .D(n29446), .Q(grid[149]) );
  LATCH grid_reg_23__4_ ( .CLK(n22505), .D(n29454), .Q(grid[142]) );
  LATCH grid_reg_23__5_ ( .CLK(n22505), .D(n29445), .Q(grid[143]) );
  LATCH grid_reg_22__4_ ( .CLK(n22502), .D(n29454), .Q(grid[136]) );
  LATCH grid_reg_22__5_ ( .CLK(n22502), .D(n29445), .Q(grid[137]) );
  LATCH grid_reg_21__4_ ( .CLK(n22499), .D(n29454), .Q(grid[130]) );
  LATCH grid_reg_21__5_ ( .CLK(n22499), .D(n29445), .Q(grid[131]) );
  LATCH grid_reg_20__4_ ( .CLK(n22496), .D(n29454), .Q(grid[124]) );
  LATCH grid_reg_20__5_ ( .CLK(n22496), .D(n29445), .Q(grid[125]) );
  LATCH grid_reg_19__4_ ( .CLK(n22493), .D(n29454), .Q(grid[118]) );
  LATCH grid_reg_19__5_ ( .CLK(n22493), .D(n29445), .Q(grid[119]) );
  LATCH grid_reg_18__4_ ( .CLK(n22490), .D(n29454), .Q(grid[112]) );
  LATCH grid_reg_18__5_ ( .CLK(n22490), .D(n29445), .Q(grid[113]) );
  LATCH grid_reg_17__4_ ( .CLK(n22487), .D(n29454), .Q(grid[106]) );
  LATCH grid_reg_17__5_ ( .CLK(n22487), .D(n29445), .Q(grid[107]) );
  LATCH grid_reg_16__4_ ( .CLK(n22484), .D(n29454), .Q(grid[100]) );
  LATCH grid_reg_16__5_ ( .CLK(n22484), .D(n29445), .Q(grid[101]) );
  LATCH grid_reg_15__4_ ( .CLK(n22481), .D(n29454), .Q(grid[94]) );
  LATCH grid_reg_15__5_ ( .CLK(n22481), .D(n29445), .Q(grid[95]) );
  LATCH grid_reg_14__4_ ( .CLK(n22478), .D(n29454), .Q(grid[88]) );
  LATCH grid_reg_14__5_ ( .CLK(n22478), .D(n29445), .Q(grid[89]) );
  LATCH grid_reg_13__4_ ( .CLK(n22475), .D(n29454), .Q(grid[82]) );
  LATCH grid_reg_13__5_ ( .CLK(n22475), .D(n29445), .Q(grid[83]) );
  LATCH grid_reg_12__4_ ( .CLK(n22472), .D(n29454), .Q(grid[76]) );
  LATCH grid_reg_12__5_ ( .CLK(n22472), .D(n29445), .Q(grid[77]) );
  LATCH grid_reg_11__4_ ( .CLK(n22469), .D(n29453), .Q(grid[70]) );
  LATCH grid_reg_11__5_ ( .CLK(n22469), .D(n29444), .Q(grid[71]) );
  LATCH grid_reg_10__4_ ( .CLK(n22466), .D(n29453), .Q(grid[64]) );
  LATCH grid_reg_10__5_ ( .CLK(n22466), .D(n29444), .Q(grid[65]) );
  LATCH grid_reg_9__4_ ( .CLK(n22463), .D(n29453), .Q(grid[58]) );
  LATCH grid_reg_9__5_ ( .CLK(n22463), .D(n29444), .Q(grid[59]) );
  LATCH grid_reg_8__4_ ( .CLK(n22460), .D(n29453), .Q(grid[52]) );
  LATCH grid_reg_8__5_ ( .CLK(n22460), .D(n29444), .Q(grid[53]) );
  LATCH grid_reg_7__4_ ( .CLK(n22457), .D(n29453), .Q(grid[46]) );
  LATCH grid_reg_7__5_ ( .CLK(n22457), .D(n29444), .Q(grid[47]) );
  LATCH grid_reg_6__4_ ( .CLK(n22454), .D(n29453), .Q(grid[40]) );
  LATCH grid_reg_6__5_ ( .CLK(n22454), .D(n29444), .Q(grid[41]) );
  LATCH grid_reg_5__4_ ( .CLK(n22451), .D(n29453), .Q(grid[34]) );
  LATCH grid_reg_5__5_ ( .CLK(n22451), .D(n29444), .Q(grid[35]) );
  LATCH grid_reg_4__4_ ( .CLK(n22448), .D(n29453), .Q(grid[28]) );
  LATCH grid_reg_4__5_ ( .CLK(n22448), .D(n29444), .Q(grid[29]) );
  LATCH grid_reg_3__4_ ( .CLK(n22445), .D(n29453), .Q(grid[22]) );
  LATCH grid_reg_3__5_ ( .CLK(n22445), .D(n29444), .Q(grid[23]) );
  LATCH grid_reg_2__4_ ( .CLK(n22442), .D(n29453), .Q(grid[16]) );
  LATCH grid_reg_2__5_ ( .CLK(n22442), .D(n29444), .Q(grid[17]) );
  LATCH grid_reg_1__4_ ( .CLK(n22439), .D(n29453), .Q(grid[10]) );
  LATCH grid_reg_1__5_ ( .CLK(n22439), .D(n29444), .Q(grid[11]) );
  LATCH grid_reg_0__4_ ( .CLK(n22436), .D(n29453), .Q(grid[4]) );
  LATCH grid_reg_0__5_ ( .CLK(n22436), .D(n29444), .Q(grid[5]) );
  LATCH addrLock_reg ( .CLK(n22429), .D(n21852), .Q(addrLock) );
  LATCH address_reg_0_ ( .CLK(n22325), .D(n21313), .Q(address[0]) );
  LATCH address_reg_1_ ( .CLK(n22325), .D(n21246), .Q(address[1]) );
  LATCH address_reg_2_ ( .CLK(n22325), .D(n21245), .Q(address[2]) );
  LATCH address_reg_3_ ( .CLK(n22325), .D(n21244), .Q(address[3]) );
  LATCH address_reg_4_ ( .CLK(n22325), .D(n21243), .Q(address[4]) );
  LATCH address_reg_5_ ( .CLK(n22325), .D(n21242), .Q(address[5]) );
  LATCH address_reg_7_ ( .CLK(n22325), .D(n29435), .Q(address[7]) );
  LATCH grid_reg_63__3_ ( .CLK(n22624), .D(n34554), .Q(grid[381]) );
  LATCH grid_reg_62__3_ ( .CLK(n22621), .D(n34553), .Q(grid[375]) );
  LATCH grid_reg_61__3_ ( .CLK(n22618), .D(n34552), .Q(grid[369]) );
  LATCH grid_reg_60__3_ ( .CLK(n22615), .D(n34551), .Q(grid[363]) );
  LATCH grid_reg_59__3_ ( .CLK(n22612), .D(n34550), .Q(grid[357]) );
  LATCH grid_reg_58__3_ ( .CLK(n22609), .D(n34549), .Q(grid[351]) );
  LATCH grid_reg_57__3_ ( .CLK(n22606), .D(n34548), .Q(grid[345]) );
  LATCH grid_reg_56__3_ ( .CLK(n22603), .D(n34547), .Q(grid[339]) );
  LATCH grid_reg_55__3_ ( .CLK(n22600), .D(n34546), .Q(grid[333]) );
  LATCH grid_reg_54__3_ ( .CLK(n22597), .D(n34545), .Q(grid[327]) );
  LATCH grid_reg_53__3_ ( .CLK(n22594), .D(n34544), .Q(grid[321]) );
  LATCH grid_reg_52__3_ ( .CLK(n22591), .D(n34543), .Q(grid[315]) );
  LATCH grid_reg_51__3_ ( .CLK(n22588), .D(n34542), .Q(grid[309]) );
  LATCH grid_reg_50__3_ ( .CLK(n22585), .D(n34541), .Q(grid[303]) );
  LATCH grid_reg_49__3_ ( .CLK(n22582), .D(n34540), .Q(grid[297]) );
  LATCH grid_reg_48__3_ ( .CLK(n22579), .D(n34539), .Q(grid[291]) );
  LATCH grid_reg_47__3_ ( .CLK(n22576), .D(n34538), .Q(grid[285]) );
  LATCH grid_reg_46__3_ ( .CLK(n22573), .D(n22242), .Q(grid[279]) );
  LATCH grid_reg_45__3_ ( .CLK(n22570), .D(n34537), .Q(grid[273]) );
  LATCH grid_reg_44__3_ ( .CLK(n22567), .D(n22234), .Q(grid[267]) );
  LATCH grid_reg_43__3_ ( .CLK(n22564), .D(n34536), .Q(grid[261]) );
  LATCH grid_reg_42__3_ ( .CLK(n22561), .D(n22226), .Q(grid[255]) );
  LATCH grid_reg_41__3_ ( .CLK(n22558), .D(n34535), .Q(grid[249]) );
  LATCH grid_reg_40__3_ ( .CLK(n22555), .D(n22218), .Q(grid[243]) );
  LATCH grid_reg_39__3_ ( .CLK(n22552), .D(n34534), .Q(grid[237]) );
  LATCH grid_reg_38__3_ ( .CLK(n22549), .D(n22210), .Q(grid[231]) );
  LATCH grid_reg_37__3_ ( .CLK(n22546), .D(n34533), .Q(grid[225]) );
  LATCH grid_reg_36__3_ ( .CLK(n22543), .D(n22202), .Q(grid[219]) );
  LATCH grid_reg_35__3_ ( .CLK(n22540), .D(n34532), .Q(grid[213]) );
  LATCH grid_reg_34__3_ ( .CLK(n22537), .D(n22194), .Q(grid[207]) );
  LATCH grid_reg_33__3_ ( .CLK(n22534), .D(n34531), .Q(grid[201]) );
  LATCH grid_reg_32__3_ ( .CLK(n22531), .D(n22186), .Q(grid[195]) );
  LATCH grid_reg_31__3_ ( .CLK(n22528), .D(n34530), .Q(grid[189]) );
  LATCH grid_reg_30__3_ ( .CLK(n22525), .D(n34529), .Q(grid[183]) );
  LATCH grid_reg_29__3_ ( .CLK(n22522), .D(n34528), .Q(grid[177]) );
  LATCH grid_reg_28__3_ ( .CLK(n22519), .D(n34527), .Q(grid[171]) );
  LATCH grid_reg_27__3_ ( .CLK(n22516), .D(n34526), .Q(grid[165]) );
  LATCH grid_reg_26__3_ ( .CLK(n22513), .D(n34525), .Q(grid[159]) );
  LATCH grid_reg_25__3_ ( .CLK(n22510), .D(n34524), .Q(grid[153]) );
  LATCH grid_reg_24__3_ ( .CLK(n22507), .D(n34523), .Q(grid[147]) );
  LATCH grid_reg_23__3_ ( .CLK(n22504), .D(n34522), .Q(grid[141]) );
  LATCH grid_reg_22__3_ ( .CLK(n22501), .D(n34521), .Q(grid[135]) );
  LATCH grid_reg_21__3_ ( .CLK(n22498), .D(n34520), .Q(grid[129]) );
  LATCH grid_reg_20__3_ ( .CLK(n22495), .D(n34519), .Q(grid[123]) );
  LATCH grid_reg_19__3_ ( .CLK(n22492), .D(n34518), .Q(grid[117]) );
  LATCH grid_reg_18__3_ ( .CLK(n22489), .D(n34517), .Q(grid[111]) );
  LATCH grid_reg_17__3_ ( .CLK(n22486), .D(n34516), .Q(grid[105]) );
  LATCH grid_reg_16__3_ ( .CLK(n22483), .D(n34515), .Q(grid[99]) );
  LATCH grid_reg_15__3_ ( .CLK(n22480), .D(n34514), .Q(grid[93]) );
  LATCH grid_reg_14__3_ ( .CLK(n22477), .D(n22114), .Q(grid[87]) );
  LATCH grid_reg_13__3_ ( .CLK(n22474), .D(n34513), .Q(grid[81]) );
  LATCH grid_reg_12__3_ ( .CLK(n22471), .D(n22106), .Q(grid[75]) );
  LATCH grid_reg_11__3_ ( .CLK(n22468), .D(n34512), .Q(grid[69]) );
  LATCH grid_reg_10__3_ ( .CLK(n22465), .D(n22098), .Q(grid[63]) );
  LATCH grid_reg_9__3_ ( .CLK(n22462), .D(n34511), .Q(grid[57]) );
  LATCH grid_reg_8__3_ ( .CLK(n22459), .D(n22090), .Q(grid[51]) );
  LATCH grid_reg_7__3_ ( .CLK(n22456), .D(n34510), .Q(grid[45]) );
  LATCH grid_reg_6__3_ ( .CLK(n22453), .D(n22082), .Q(grid[39]) );
  LATCH grid_reg_5__3_ ( .CLK(n22450), .D(n34509), .Q(grid[33]) );
  LATCH grid_reg_4__3_ ( .CLK(n22447), .D(n22074), .Q(grid[27]) );
  LATCH grid_reg_3__3_ ( .CLK(n22444), .D(n34508), .Q(grid[21]) );
  LATCH grid_reg_2__3_ ( .CLK(n22441), .D(n22066), .Q(grid[15]) );
  LATCH grid_reg_1__3_ ( .CLK(n22438), .D(n34507), .Q(grid[9]) );
  LATCH grid_reg_0__3_ ( .CLK(n22435), .D(n22056), .Q(grid[3]) );
  LATCH grid_reg_63__0_ ( .CLK(n22624), .D(n23269), .Q(grid[378]) );
  LATCH grid_reg_63__1_ ( .CLK(n22624), .D(n22308), .Q(grid[379]) );
  LATCH grid_reg_63__2_ ( .CLK(n22624), .D(n22309), .Q(grid[380]) );
  LATCH grid_reg_62__0_ ( .CLK(n22621), .D(n22303), .Q(grid[372]) );
  LATCH grid_reg_62__1_ ( .CLK(n22621), .D(n22304), .Q(grid[373]) );
  LATCH grid_reg_62__2_ ( .CLK(n22621), .D(n22305), .Q(grid[374]) );
  LATCH grid_reg_61__0_ ( .CLK(n22618), .D(n22299), .Q(grid[366]) );
  LATCH grid_reg_61__1_ ( .CLK(n22618), .D(n22300), .Q(grid[367]) );
  LATCH grid_reg_61__2_ ( .CLK(n22618), .D(n22301), .Q(grid[368]) );
  LATCH grid_reg_60__0_ ( .CLK(n22615), .D(n22295), .Q(grid[360]) );
  LATCH grid_reg_60__1_ ( .CLK(n22615), .D(n22296), .Q(grid[361]) );
  LATCH grid_reg_60__2_ ( .CLK(n22615), .D(n22297), .Q(grid[362]) );
  LATCH grid_reg_59__0_ ( .CLK(n22612), .D(n22291), .Q(grid[354]) );
  LATCH grid_reg_59__1_ ( .CLK(n22612), .D(n22292), .Q(grid[355]) );
  LATCH grid_reg_59__2_ ( .CLK(n22612), .D(n22293), .Q(grid[356]) );
  LATCH grid_reg_58__0_ ( .CLK(n22609), .D(n22287), .Q(grid[348]) );
  LATCH grid_reg_58__1_ ( .CLK(n22609), .D(n22288), .Q(grid[349]) );
  LATCH grid_reg_58__2_ ( .CLK(n22609), .D(n22289), .Q(grid[350]) );
  LATCH grid_reg_57__0_ ( .CLK(n22606), .D(n22283), .Q(grid[342]) );
  LATCH grid_reg_57__1_ ( .CLK(n22606), .D(n22284), .Q(grid[343]) );
  LATCH grid_reg_57__2_ ( .CLK(n22606), .D(n22285), .Q(grid[344]) );
  LATCH grid_reg_56__0_ ( .CLK(n22603), .D(n22279), .Q(grid[336]) );
  LATCH grid_reg_56__1_ ( .CLK(n22603), .D(n22280), .Q(grid[337]) );
  LATCH grid_reg_56__2_ ( .CLK(n22603), .D(n22281), .Q(grid[338]) );
  LATCH grid_reg_55__0_ ( .CLK(n22600), .D(n22275), .Q(grid[330]) );
  LATCH grid_reg_55__1_ ( .CLK(n22600), .D(n22276), .Q(grid[331]) );
  LATCH grid_reg_55__2_ ( .CLK(n22600), .D(n22277), .Q(grid[332]) );
  LATCH grid_reg_54__0_ ( .CLK(n22597), .D(n22271), .Q(grid[324]) );
  LATCH grid_reg_54__1_ ( .CLK(n22597), .D(n22272), .Q(grid[325]) );
  LATCH grid_reg_54__2_ ( .CLK(n22597), .D(n23266), .Q(grid[326]) );
  LATCH grid_reg_53__0_ ( .CLK(n22594), .D(n22267), .Q(grid[318]) );
  LATCH grid_reg_53__1_ ( .CLK(n22594), .D(n22268), .Q(grid[319]) );
  LATCH grid_reg_53__2_ ( .CLK(n22594), .D(n22269), .Q(grid[320]) );
  LATCH grid_reg_52__0_ ( .CLK(n22591), .D(n22263), .Q(grid[312]) );
  LATCH grid_reg_52__1_ ( .CLK(n22591), .D(n22264), .Q(grid[313]) );
  LATCH grid_reg_52__2_ ( .CLK(n22591), .D(n23262), .Q(grid[314]) );
  LATCH grid_reg_51__0_ ( .CLK(n22588), .D(n22259), .Q(grid[306]) );
  LATCH grid_reg_51__1_ ( .CLK(n22588), .D(n22260), .Q(grid[307]) );
  LATCH grid_reg_51__2_ ( .CLK(n22588), .D(n22261), .Q(grid[308]) );
  LATCH grid_reg_50__0_ ( .CLK(n22585), .D(n22255), .Q(grid[300]) );
  LATCH grid_reg_50__1_ ( .CLK(n22585), .D(n22256), .Q(grid[301]) );
  LATCH grid_reg_50__2_ ( .CLK(n22585), .D(n22257), .Q(grid[302]) );
  LATCH grid_reg_49__0_ ( .CLK(n22582), .D(n22251), .Q(grid[294]) );
  LATCH grid_reg_49__1_ ( .CLK(n22582), .D(n22252), .Q(grid[295]) );
  LATCH grid_reg_49__2_ ( .CLK(n22582), .D(n22253), .Q(grid[296]) );
  LATCH grid_reg_48__0_ ( .CLK(n22579), .D(n22247), .Q(grid[288]) );
  LATCH grid_reg_48__1_ ( .CLK(n22579), .D(n22248), .Q(grid[289]) );
  LATCH grid_reg_48__2_ ( .CLK(n22579), .D(n22249), .Q(grid[290]) );
  LATCH grid_reg_47__0_ ( .CLK(n22576), .D(n22243), .Q(grid[282]) );
  LATCH grid_reg_47__1_ ( .CLK(n22576), .D(n22244), .Q(grid[283]) );
  LATCH grid_reg_47__2_ ( .CLK(n22576), .D(n23623), .Q(grid[284]) );
  LATCH grid_reg_46__0_ ( .CLK(n22573), .D(n22239), .Q(grid[276]) );
  LATCH grid_reg_46__1_ ( .CLK(n22573), .D(n22240), .Q(grid[277]) );
  LATCH grid_reg_46__2_ ( .CLK(n22573), .D(n23259), .Q(grid[278]) );
  LATCH grid_reg_45__0_ ( .CLK(n22570), .D(n22235), .Q(grid[270]) );
  LATCH grid_reg_45__1_ ( .CLK(n22570), .D(n22236), .Q(grid[271]) );
  LATCH grid_reg_45__2_ ( .CLK(n22570), .D(n23255), .Q(grid[272]) );
  LATCH grid_reg_44__0_ ( .CLK(n22567), .D(n22231), .Q(grid[264]) );
  LATCH grid_reg_44__1_ ( .CLK(n22567), .D(n22232), .Q(grid[265]) );
  LATCH grid_reg_44__2_ ( .CLK(n22567), .D(n22233), .Q(grid[266]) );
  LATCH grid_reg_43__0_ ( .CLK(n22564), .D(n22227), .Q(grid[258]) );
  LATCH grid_reg_43__1_ ( .CLK(n22564), .D(n22228), .Q(grid[259]) );
  LATCH grid_reg_43__2_ ( .CLK(n22564), .D(n23252), .Q(grid[260]) );
  LATCH grid_reg_42__0_ ( .CLK(n22561), .D(n22223), .Q(grid[252]) );
  LATCH grid_reg_42__1_ ( .CLK(n22561), .D(n22224), .Q(grid[253]) );
  LATCH grid_reg_42__2_ ( .CLK(n22561), .D(n22225), .Q(grid[254]) );
  LATCH grid_reg_41__0_ ( .CLK(n22558), .D(n22219), .Q(grid[246]) );
  LATCH grid_reg_41__1_ ( .CLK(n22558), .D(n22220), .Q(grid[247]) );
  LATCH grid_reg_41__2_ ( .CLK(n22558), .D(n22221), .Q(grid[248]) );
  LATCH grid_reg_40__0_ ( .CLK(n22555), .D(n22215), .Q(grid[240]) );
  LATCH grid_reg_40__1_ ( .CLK(n22555), .D(n22216), .Q(grid[241]) );
  LATCH grid_reg_40__2_ ( .CLK(n22555), .D(n22217), .Q(grid[242]) );
  LATCH grid_reg_39__0_ ( .CLK(n22552), .D(n22211), .Q(grid[234]) );
  LATCH grid_reg_39__1_ ( .CLK(n22552), .D(n22212), .Q(grid[235]) );
  LATCH grid_reg_39__2_ ( .CLK(n22552), .D(n22213), .Q(grid[236]) );
  LATCH grid_reg_38__0_ ( .CLK(n22549), .D(n22207), .Q(grid[228]) );
  LATCH grid_reg_38__1_ ( .CLK(n22549), .D(n22208), .Q(grid[229]) );
  LATCH grid_reg_38__2_ ( .CLK(n22549), .D(n22209), .Q(grid[230]) );
  LATCH grid_reg_37__0_ ( .CLK(n22546), .D(n22203), .Q(grid[222]) );
  LATCH grid_reg_37__1_ ( .CLK(n22546), .D(n22204), .Q(grid[223]) );
  LATCH grid_reg_37__2_ ( .CLK(n22546), .D(n22205), .Q(grid[224]) );
  LATCH grid_reg_36__0_ ( .CLK(n22543), .D(n22199), .Q(grid[216]) );
  LATCH grid_reg_36__1_ ( .CLK(n22543), .D(n22200), .Q(grid[217]) );
  LATCH grid_reg_36__2_ ( .CLK(n22543), .D(n22201), .Q(grid[218]) );
  LATCH grid_reg_35__0_ ( .CLK(n22540), .D(n22195), .Q(grid[210]) );
  LATCH grid_reg_35__1_ ( .CLK(n22540), .D(n22196), .Q(grid[211]) );
  LATCH grid_reg_35__2_ ( .CLK(n22540), .D(n22197), .Q(grid[212]) );
  LATCH grid_reg_34__0_ ( .CLK(n22537), .D(n22191), .Q(grid[204]) );
  LATCH grid_reg_34__1_ ( .CLK(n22537), .D(n22192), .Q(grid[205]) );
  LATCH grid_reg_34__2_ ( .CLK(n22537), .D(n22193), .Q(grid[206]) );
  LATCH grid_reg_33__0_ ( .CLK(n22534), .D(n22187), .Q(grid[198]) );
  LATCH grid_reg_33__1_ ( .CLK(n22534), .D(n22188), .Q(grid[199]) );
  LATCH grid_reg_33__2_ ( .CLK(n22534), .D(n22189), .Q(grid[200]) );
  LATCH grid_reg_32__0_ ( .CLK(n22531), .D(n22183), .Q(grid[192]) );
  LATCH grid_reg_32__1_ ( .CLK(n22531), .D(n22184), .Q(grid[193]) );
  LATCH grid_reg_32__2_ ( .CLK(n22531), .D(n22185), .Q(grid[194]) );
  LATCH grid_reg_31__0_ ( .CLK(n22528), .D(n22179), .Q(grid[186]) );
  LATCH grid_reg_31__1_ ( .CLK(n22528), .D(n22180), .Q(grid[187]) );
  LATCH grid_reg_31__2_ ( .CLK(n22528), .D(n22181), .Q(grid[188]) );
  LATCH grid_reg_30__0_ ( .CLK(n22525), .D(n22175), .Q(grid[180]) );
  LATCH grid_reg_30__1_ ( .CLK(n22525), .D(n22176), .Q(grid[181]) );
  LATCH grid_reg_30__2_ ( .CLK(n22525), .D(n23249), .Q(grid[182]) );
  LATCH grid_reg_29__0_ ( .CLK(n22522), .D(n22171), .Q(grid[174]) );
  LATCH grid_reg_29__1_ ( .CLK(n22522), .D(n22172), .Q(grid[175]) );
  LATCH grid_reg_29__2_ ( .CLK(n22522), .D(n22173), .Q(grid[176]) );
  LATCH grid_reg_28__0_ ( .CLK(n22519), .D(n22167), .Q(grid[168]) );
  LATCH grid_reg_28__1_ ( .CLK(n22519), .D(n22168), .Q(grid[169]) );
  LATCH grid_reg_28__2_ ( .CLK(n22519), .D(n23246), .Q(grid[170]) );
  LATCH grid_reg_27__0_ ( .CLK(n22516), .D(n22163), .Q(grid[162]) );
  LATCH grid_reg_27__1_ ( .CLK(n22516), .D(n22164), .Q(grid[163]) );
  LATCH grid_reg_27__2_ ( .CLK(n22516), .D(n22165), .Q(grid[164]) );
  LATCH grid_reg_26__0_ ( .CLK(n22513), .D(n22159), .Q(grid[156]) );
  LATCH grid_reg_26__1_ ( .CLK(n22513), .D(n22160), .Q(grid[157]) );
  LATCH grid_reg_26__2_ ( .CLK(n22513), .D(n22161), .Q(grid[158]) );
  LATCH grid_reg_25__0_ ( .CLK(n22510), .D(n22155), .Q(grid[150]) );
  LATCH grid_reg_25__1_ ( .CLK(n22510), .D(n22156), .Q(grid[151]) );
  LATCH grid_reg_25__2_ ( .CLK(n22510), .D(n22157), .Q(grid[152]) );
  LATCH grid_reg_24__0_ ( .CLK(n22507), .D(n22151), .Q(grid[144]) );
  LATCH grid_reg_24__1_ ( .CLK(n22507), .D(n22152), .Q(grid[145]) );
  LATCH grid_reg_24__2_ ( .CLK(n22507), .D(n22153), .Q(grid[146]) );
  LATCH grid_reg_23__0_ ( .CLK(n22504), .D(n22147), .Q(grid[138]) );
  LATCH grid_reg_23__1_ ( .CLK(n22504), .D(n22148), .Q(grid[139]) );
  LATCH grid_reg_23__2_ ( .CLK(n22504), .D(n22149), .Q(grid[140]) );
  LATCH grid_reg_22__0_ ( .CLK(n22501), .D(n22143), .Q(grid[132]) );
  LATCH grid_reg_22__1_ ( .CLK(n22501), .D(n22144), .Q(grid[133]) );
  LATCH grid_reg_22__2_ ( .CLK(n22501), .D(n23243), .Q(grid[134]) );
  LATCH grid_reg_21__0_ ( .CLK(n22498), .D(n22139), .Q(grid[126]) );
  LATCH grid_reg_21__1_ ( .CLK(n22498), .D(n22140), .Q(grid[127]) );
  LATCH grid_reg_21__2_ ( .CLK(n22498), .D(n22141), .Q(grid[128]) );
  LATCH grid_reg_20__0_ ( .CLK(n22495), .D(n22135), .Q(grid[120]) );
  LATCH grid_reg_20__1_ ( .CLK(n22495), .D(n22136), .Q(grid[121]) );
  LATCH grid_reg_20__2_ ( .CLK(n22495), .D(n22137), .Q(grid[122]) );
  LATCH grid_reg_19__0_ ( .CLK(n22492), .D(n22131), .Q(grid[114]) );
  LATCH grid_reg_19__1_ ( .CLK(n22492), .D(n22132), .Q(grid[115]) );
  LATCH grid_reg_19__2_ ( .CLK(n22492), .D(n22133), .Q(grid[116]) );
  LATCH grid_reg_18__0_ ( .CLK(n22489), .D(n22127), .Q(grid[108]) );
  LATCH grid_reg_18__1_ ( .CLK(n22489), .D(n22128), .Q(grid[109]) );
  LATCH grid_reg_18__2_ ( .CLK(n22489), .D(n23620), .Q(grid[110]) );
  LATCH grid_reg_17__0_ ( .CLK(n22486), .D(n22123), .Q(grid[102]) );
  LATCH grid_reg_17__1_ ( .CLK(n22486), .D(n22124), .Q(grid[103]) );
  LATCH grid_reg_17__2_ ( .CLK(n22486), .D(n22125), .Q(grid[104]) );
  LATCH grid_reg_16__0_ ( .CLK(n22483), .D(n22119), .Q(grid[96]) );
  LATCH grid_reg_16__1_ ( .CLK(n22483), .D(n22120), .Q(grid[97]) );
  LATCH grid_reg_16__2_ ( .CLK(n22483), .D(n22121), .Q(grid[98]) );
  LATCH grid_reg_15__0_ ( .CLK(n22480), .D(n22115), .Q(grid[90]) );
  LATCH grid_reg_15__1_ ( .CLK(n22480), .D(n22116), .Q(grid[91]) );
  LATCH grid_reg_15__2_ ( .CLK(n22480), .D(n22117), .Q(grid[92]) );
  LATCH grid_reg_14__0_ ( .CLK(n22477), .D(n22111), .Q(grid[84]) );
  LATCH grid_reg_14__1_ ( .CLK(n22477), .D(n22112), .Q(grid[85]) );
  LATCH grid_reg_14__2_ ( .CLK(n22477), .D(n23617), .Q(grid[86]) );
  LATCH grid_reg_13__0_ ( .CLK(n22474), .D(n22107), .Q(grid[78]) );
  LATCH grid_reg_13__1_ ( .CLK(n22474), .D(n22108), .Q(grid[79]) );
  LATCH grid_reg_13__2_ ( .CLK(n22474), .D(n23240), .Q(grid[80]) );
  LATCH grid_reg_12__0_ ( .CLK(n22471), .D(n22103), .Q(grid[72]) );
  LATCH grid_reg_12__1_ ( .CLK(n22471), .D(n22104), .Q(grid[73]) );
  LATCH grid_reg_12__2_ ( .CLK(n22471), .D(n22105), .Q(grid[74]) );
  LATCH grid_reg_11__0_ ( .CLK(n22468), .D(n22099), .Q(grid[66]) );
  LATCH grid_reg_11__1_ ( .CLK(n22468), .D(n22100), .Q(grid[67]) );
  LATCH grid_reg_11__2_ ( .CLK(n22468), .D(n22101), .Q(grid[68]) );
  LATCH grid_reg_10__0_ ( .CLK(n22465), .D(n22095), .Q(grid[60]) );
  LATCH grid_reg_10__1_ ( .CLK(n22465), .D(n22096), .Q(grid[61]) );
  LATCH grid_reg_10__2_ ( .CLK(n22465), .D(n23237), .Q(grid[62]) );
  LATCH grid_reg_9__0_ ( .CLK(n22462), .D(n22091), .Q(grid[54]) );
  LATCH grid_reg_9__1_ ( .CLK(n22462), .D(n22092), .Q(grid[55]) );
  LATCH grid_reg_9__2_ ( .CLK(n22462), .D(n22093), .Q(grid[56]) );
  LATCH grid_reg_8__0_ ( .CLK(n22459), .D(n22087), .Q(grid[48]) );
  LATCH grid_reg_8__1_ ( .CLK(n22459), .D(n22088), .Q(grid[49]) );
  LATCH grid_reg_8__2_ ( .CLK(n22459), .D(n23234), .Q(grid[50]) );
  LATCH grid_reg_7__0_ ( .CLK(n22456), .D(n22083), .Q(grid[42]) );
  LATCH grid_reg_7__1_ ( .CLK(n22456), .D(n22084), .Q(grid[43]) );
  LATCH grid_reg_7__2_ ( .CLK(n22456), .D(n23230), .Q(grid[44]) );
  LATCH grid_reg_6__0_ ( .CLK(n22453), .D(n22079), .Q(grid[36]) );
  LATCH grid_reg_6__1_ ( .CLK(n22453), .D(n22080), .Q(grid[37]) );
  LATCH grid_reg_6__2_ ( .CLK(n22453), .D(n23227), .Q(grid[38]) );
  LATCH grid_reg_5__0_ ( .CLK(n22450), .D(n22075), .Q(grid[30]) );
  LATCH grid_reg_5__1_ ( .CLK(n22450), .D(n22076), .Q(grid[31]) );
  LATCH grid_reg_5__2_ ( .CLK(n22450), .D(n23223), .Q(grid[32]) );
  LATCH grid_reg_4__0_ ( .CLK(n22447), .D(n22071), .Q(grid[24]) );
  LATCH grid_reg_4__1_ ( .CLK(n22447), .D(n22072), .Q(grid[25]) );
  LATCH grid_reg_4__2_ ( .CLK(n22447), .D(n23220), .Q(grid[26]) );
  LATCH grid_reg_3__0_ ( .CLK(n22444), .D(n22067), .Q(grid[18]) );
  LATCH grid_reg_3__1_ ( .CLK(n22444), .D(n22068), .Q(grid[19]) );
  LATCH grid_reg_3__2_ ( .CLK(n22444), .D(n23217), .Q(grid[20]) );
  LATCH grid_reg_2__0_ ( .CLK(n22441), .D(n22063), .Q(grid[12]) );
  LATCH grid_reg_2__1_ ( .CLK(n22441), .D(n22064), .Q(grid[13]) );
  LATCH grid_reg_2__2_ ( .CLK(n22441), .D(n23214), .Q(grid[14]) );
  LATCH grid_reg_1__0_ ( .CLK(n22438), .D(n22059), .Q(grid[6]) );
  LATCH grid_reg_1__1_ ( .CLK(n22438), .D(n22060), .Q(grid[7]) );
  LATCH grid_reg_1__2_ ( .CLK(n22438), .D(n23211), .Q(grid[8]) );
  LATCH grid_reg_0__0_ ( .CLK(n22435), .D(n22053), .Q(grid[0]) );
  LATCH grid_reg_0__1_ ( .CLK(n22435), .D(n22054), .Q(grid[1]) );
  LATCH grid_reg_0__2_ ( .CLK(n22435), .D(n22055), .Q(grid[2]) );
  AND2X2 U19 ( .A(n34555), .B(n22635), .Y(n22634) );
  AND2X2 U20 ( .A(n27304), .B(n22635), .Y(n22633) );
  AND2X2 U22 ( .A(n25466), .B(n14097), .Y(n22635) );
  AND2X2 U86 ( .A(n29220), .B(n15155), .Y(n14369) );
  AND2X2 U87 ( .A(n15155), .B(n34498), .Y(n14368) );
  AND2X2 U89 ( .A(n29440), .B(n14097), .Y(n14371) );
  AND2X2 U94 ( .A(n26895), .B(n2219), .Y(n15183) );
  AND2X2 U95 ( .A(n15155), .B(n20818), .Y(n15182) );
  AND2X2 U96 ( .A(net64168), .B(n14097), .Y(n15155) );
  OR2X2 U97 ( .A(n15226), .B(n14218), .Y(n22419) );
  OR2X2 U99 ( .A(n15235), .B(n14218), .Y(n22418) );
  OR2X2 U101 ( .A(n15256), .B(n14218), .Y(n22416) );
  OR2X2 U102 ( .A(n15279), .B(n14218), .Y(n22413) );
  OR2X2 U103 ( .A(n15302), .B(n14218), .Y(n22410) );
  OR2X2 U104 ( .A(n15325), .B(n14218), .Y(n22407) );
  OR2X2 U105 ( .A(n15348), .B(n14218), .Y(n22404) );
  OR2X2 U107 ( .A(n15373), .B(n14218), .Y(n22401) );
  OR2X2 U108 ( .A(n15397), .B(n14218), .Y(n22398) );
  OR2X2 U109 ( .A(n15420), .B(n14218), .Y(n22395) );
  OR2X2 U110 ( .A(n15442), .B(n14218), .Y(n22392) );
  OR2X2 U111 ( .A(n15464), .B(n14218), .Y(n22389) );
  OR2X2 U112 ( .A(n15486), .B(n14218), .Y(n22386) );
  OR2X2 U113 ( .A(n15508), .B(n14218), .Y(n22383) );
  OR2X2 U114 ( .A(n15529), .B(n14218), .Y(n22380) );
  OR2X2 U120 ( .A(n15597), .B(n14218), .Y(n22370) );
  OR2X2 U121 ( .A(n15618), .B(n14218), .Y(n22367) );
  OR2X2 U122 ( .A(n15639), .B(n14218), .Y(n22364) );
  OR2X2 U123 ( .A(n15660), .B(n14218), .Y(n22361) );
  OR2X2 U124 ( .A(n15681), .B(n14218), .Y(n22358) );
  OR2X2 U125 ( .A(n15702), .B(n14218), .Y(n22355) );
  OR2X2 U127 ( .A(n15724), .B(n14218), .Y(n22352) );
  OR2X2 U128 ( .A(n15746), .B(n14218), .Y(n22349) );
  OR2X2 U129 ( .A(n15767), .B(n14218), .Y(n22346) );
  OR2X2 U130 ( .A(n15788), .B(n14218), .Y(n22343) );
  OR2X2 U131 ( .A(n15809), .B(n14218), .Y(n22340) );
  OR2X2 U132 ( .A(n15830), .B(n14218), .Y(n22337) );
  OR2X2 U133 ( .A(n15851), .B(n14218), .Y(n22334) );
  INVX2 U288 ( .A(clk), .Y(n2219) );
  INVX2 U1897 ( .A(n14373), .Y(n14097) );
  INVX2 U2018 ( .A(n15201), .Y(n14218) );
  NAND3X1 U2140 ( .A(n13743), .B(n14349), .C(n14350), .Y(n22632) );
  AOI22X1 U2141 ( .A(n14351), .B(n23281), .C(n34498), .D(n22635), .Y(n14350)
         );
  NOR3X1 U2142 ( .A(n14346), .B(n14348), .C(n24922), .Y(n14354) );
  OAI21X1 U2143 ( .A(n14356), .B(net108619), .C(n14349), .Y(n22631) );
  OAI21X1 U2144 ( .A(n14356), .B(net109176), .C(n14349), .Y(n22630) );
  OAI21X1 U2145 ( .A(n14356), .B(n26062), .C(n14349), .Y(n22629) );
  OAI21X1 U2146 ( .A(n14356), .B(net110410), .C(n14349), .Y(n22628) );
  NAND2X1 U2147 ( .A(n22635), .B(n29191), .Y(n14349) );
  NAND2X1 U2148 ( .A(n20818), .B(n22635), .Y(n14356) );
  NAND2X1 U2151 ( .A(n14097), .B(net96340), .Y(n14348) );
  AOI22X1 U2153 ( .A(n34495), .B(n14368), .C(n34496), .D(n14369), .Y(n14366)
         );
  OAI21X1 U2156 ( .A(n24281), .B(n14373), .C(n14374), .Y(n22624) );
  AOI21X1 U2157 ( .A(n34603), .B(1'b0), .C(n14218), .Y(n14374) );
  NAND3X1 U2161 ( .A(n14384), .B(n34604), .C(cs), .Y(n14382) );
  OAI21X1 U2167 ( .A(n14390), .B(n14373), .C(n14391), .Y(n22621) );
  AOI21X1 U2168 ( .A(n30466), .B(1'b0), .C(n14218), .Y(n14391) );
  NAND3X1 U2172 ( .A(cs), .B(n34604), .C(n14398), .Y(n14396) );
  OAI21X1 U2178 ( .A(n14403), .B(n14373), .C(n14404), .Y(n22618) );
  AOI21X1 U2179 ( .A(n34602), .B(1'b0), .C(n14218), .Y(n14404) );
  NAND3X1 U2183 ( .A(cs), .B(n34604), .C(n14411), .Y(n14409) );
  OAI21X1 U2189 ( .A(n14416), .B(n14373), .C(n14417), .Y(n22615) );
  AOI21X1 U2190 ( .A(n30452), .B(1'b0), .C(n14218), .Y(n14417) );
  NAND3X1 U2194 ( .A(cs), .B(n34604), .C(n14424), .Y(n14422) );
  OAI21X1 U2200 ( .A(n14429), .B(n14373), .C(n14430), .Y(n22612) );
  AOI21X1 U2201 ( .A(n30444), .B(1'b0), .C(n14218), .Y(n14430) );
  NAND3X1 U2205 ( .A(cs), .B(n34604), .C(n14437), .Y(n14435) );
  OAI21X1 U2211 ( .A(n14442), .B(n14373), .C(n14443), .Y(n22609) );
  AOI21X1 U2212 ( .A(n30435), .B(1'b0), .C(n14218), .Y(n14443) );
  NAND3X1 U2216 ( .A(cs), .B(n34604), .C(n14450), .Y(n14448) );
  OAI21X1 U2222 ( .A(n14455), .B(n14373), .C(n14456), .Y(n22606) );
  AOI21X1 U2223 ( .A(n30427), .B(1'b0), .C(n14218), .Y(n14456) );
  NAND3X1 U2227 ( .A(cs), .B(n34604), .C(n14463), .Y(n14461) );
  OAI21X1 U2233 ( .A(n14468), .B(n14373), .C(n14469), .Y(n22603) );
  AOI21X1 U2234 ( .A(n30421), .B(1'b0), .C(n14218), .Y(n14469) );
  NAND3X1 U2238 ( .A(cs), .B(n34604), .C(n14476), .Y(n14474) );
  NAND3X1 U2239 ( .A(n20975), .B(n20812), .C(n26985), .Y(n14477) );
  OAI21X1 U2245 ( .A(n14483), .B(n14373), .C(n14484), .Y(n22600) );
  AOI21X1 U2246 ( .A(n30413), .B(1'b0), .C(n14218), .Y(n14484) );
  NAND3X1 U2250 ( .A(cs), .B(n14384), .C(n34600), .Y(n14489) );
  OAI21X1 U2256 ( .A(n14495), .B(n14373), .C(n14496), .Y(n22597) );
  AOI21X1 U2257 ( .A(n30404), .B(1'b0), .C(n14218), .Y(n14496) );
  NAND3X1 U2261 ( .A(n14398), .B(cs), .C(n34600), .Y(n14501) );
  OAI21X1 U2267 ( .A(n14507), .B(n14373), .C(n14508), .Y(n22594) );
  AOI21X1 U2268 ( .A(n30399), .B(1'b0), .C(n14218), .Y(n14508) );
  NAND3X1 U2272 ( .A(n14411), .B(cs), .C(n34600), .Y(n14513) );
  OAI21X1 U2278 ( .A(n14519), .B(n14373), .C(n14520), .Y(n22591) );
  AOI21X1 U2279 ( .A(n30394), .B(1'b0), .C(n14218), .Y(n14520) );
  NAND3X1 U2283 ( .A(n14424), .B(cs), .C(n34600), .Y(n14525) );
  OAI21X1 U2289 ( .A(n14531), .B(n14373), .C(n14532), .Y(n22588) );
  AOI21X1 U2290 ( .A(n30389), .B(1'b0), .C(n14218), .Y(n14532) );
  NAND3X1 U2294 ( .A(n14437), .B(cs), .C(n34600), .Y(n14537) );
  OAI21X1 U2300 ( .A(n14543), .B(n14373), .C(n14544), .Y(n22585) );
  AOI21X1 U2301 ( .A(n34599), .B(1'b0), .C(n14218), .Y(n14544) );
  NAND3X1 U2305 ( .A(n14450), .B(cs), .C(n34600), .Y(n14549) );
  OAI21X1 U2311 ( .A(n14555), .B(n14373), .C(n14556), .Y(n22582) );
  AOI21X1 U2312 ( .A(n30380), .B(1'b0), .C(n14218), .Y(n14556) );
  NAND3X1 U2316 ( .A(n14463), .B(cs), .C(n34600), .Y(n14561) );
  OAI21X1 U2322 ( .A(n14567), .B(n14373), .C(n14568), .Y(n22579) );
  AOI21X1 U2323 ( .A(n30375), .B(1'b0), .C(n14218), .Y(n14568) );
  NAND3X1 U2327 ( .A(n14476), .B(cs), .C(n34600), .Y(n14573) );
  NAND3X1 U2328 ( .A(n20975), .B(n20812), .C(n27063), .Y(n14575) );
  OAI21X1 U2334 ( .A(n14581), .B(n14373), .C(n14582), .Y(n22576) );
  AOI21X1 U2335 ( .A(n30366), .B(1'b0), .C(n14218), .Y(n14582) );
  NAND3X1 U2339 ( .A(cs), .B(n14384), .C(n34610), .Y(n14587) );
  OAI21X1 U2345 ( .A(n14593), .B(n14373), .C(n14594), .Y(n22573) );
  AOI21X1 U2346 ( .A(n30359), .B(1'b0), .C(n14218), .Y(n14594) );
  NAND3X1 U2350 ( .A(n14398), .B(cs), .C(n34610), .Y(n14599) );
  OAI21X1 U2356 ( .A(n14605), .B(n14373), .C(n14606), .Y(n22570) );
  AOI21X1 U2357 ( .A(n30354), .B(1'b0), .C(n14218), .Y(n14606) );
  NAND3X1 U2361 ( .A(n14411), .B(cs), .C(n34610), .Y(n14611) );
  OAI21X1 U2367 ( .A(n14617), .B(n14373), .C(n14618), .Y(n22567) );
  AOI21X1 U2368 ( .A(n30349), .B(1'b0), .C(n14218), .Y(n14618) );
  NAND3X1 U2372 ( .A(n14424), .B(cs), .C(n34610), .Y(n14623) );
  OAI21X1 U2378 ( .A(n14629), .B(n14373), .C(n14630), .Y(n22564) );
  AOI21X1 U2379 ( .A(n34609), .B(1'b0), .C(n14218), .Y(n14630) );
  NAND3X1 U2383 ( .A(n14437), .B(cs), .C(n34610), .Y(n14635) );
  OAI21X1 U2389 ( .A(n14641), .B(n14373), .C(n14642), .Y(n22561) );
  AOI21X1 U2390 ( .A(n30340), .B(1'b0), .C(n14218), .Y(n14642) );
  NAND3X1 U2394 ( .A(n14450), .B(cs), .C(n34610), .Y(n14647) );
  OAI21X1 U2400 ( .A(n14653), .B(n14373), .C(n14654), .Y(n22558) );
  AOI21X1 U2401 ( .A(n30335), .B(1'b0), .C(n14218), .Y(n14654) );
  NAND3X1 U2405 ( .A(n14463), .B(cs), .C(n34610), .Y(n14659) );
  OAI21X1 U2411 ( .A(n14665), .B(n14373), .C(n14666), .Y(n22555) );
  AOI21X1 U2412 ( .A(n30330), .B(1'b0), .C(n14218), .Y(n14666) );
  NAND3X1 U2416 ( .A(n14476), .B(cs), .C(n34610), .Y(n14671) );
  NAND3X1 U2417 ( .A(n20975), .B(address[3]), .C(n21402), .Y(n14673) );
  OAI21X1 U2424 ( .A(n14680), .B(n14373), .C(n14681), .Y(n22552) );
  AOI21X1 U2425 ( .A(n30322), .B(1'b0), .C(n14218), .Y(n14681) );
  NAND3X1 U2429 ( .A(cs), .B(n14384), .C(n34608), .Y(n14686) );
  OAI21X1 U2435 ( .A(n14692), .B(n14373), .C(n14693), .Y(n22549) );
  AOI21X1 U2436 ( .A(n30314), .B(1'b0), .C(n14218), .Y(n14693) );
  NAND3X1 U2440 ( .A(n14398), .B(cs), .C(n34608), .Y(n14698) );
  OAI21X1 U2446 ( .A(n14704), .B(n14373), .C(n14705), .Y(n22546) );
  AOI21X1 U2447 ( .A(n30309), .B(1'b0), .C(n14218), .Y(n14705) );
  NAND3X1 U2451 ( .A(n14411), .B(cs), .C(n34608), .Y(n14710) );
  OAI21X1 U2457 ( .A(n14716), .B(n14373), .C(n14717), .Y(n22543) );
  AOI21X1 U2458 ( .A(n30304), .B(1'b0), .C(n14218), .Y(n14717) );
  NAND3X1 U2462 ( .A(n14424), .B(cs), .C(n34608), .Y(n14722) );
  OAI21X1 U2468 ( .A(n14728), .B(n14373), .C(n14729), .Y(n22540) );
  AOI21X1 U2469 ( .A(n30299), .B(1'b0), .C(n14218), .Y(n14729) );
  NAND3X1 U2473 ( .A(n14437), .B(cs), .C(n34608), .Y(n14734) );
  OAI21X1 U2479 ( .A(n14740), .B(n14373), .C(n14741), .Y(n22537) );
  AOI21X1 U2480 ( .A(n30294), .B(1'b0), .C(n14218), .Y(n14741) );
  NAND3X1 U2484 ( .A(n14450), .B(cs), .C(n34608), .Y(n14746) );
  OAI21X1 U2490 ( .A(n14752), .B(n14373), .C(n14753), .Y(n22534) );
  AOI21X1 U2491 ( .A(n30289), .B(1'b0), .C(n14218), .Y(n14753) );
  NAND3X1 U2495 ( .A(n14463), .B(cs), .C(n34608), .Y(n14758) );
  OAI21X1 U2501 ( .A(n14764), .B(n14373), .C(n14765), .Y(n22531) );
  AOI21X1 U2502 ( .A(n30284), .B(1'b0), .C(n14218), .Y(n14765) );
  NAND3X1 U2506 ( .A(n14476), .B(cs), .C(n34608), .Y(n14770) );
  NAND3X1 U2507 ( .A(n29469), .B(n34615), .C(n24877), .Y(n14772) );
  OAI21X1 U2514 ( .A(n14778), .B(n14373), .C(n14779), .Y(n22528) );
  AOI21X1 U2515 ( .A(n30275), .B(1'b0), .C(n14218), .Y(n14779) );
  NAND3X1 U2519 ( .A(cs), .B(n14384), .C(n34607), .Y(n14784) );
  OAI21X1 U2525 ( .A(n14790), .B(n14373), .C(n14791), .Y(n22525) );
  AOI21X1 U2526 ( .A(n34606), .B(1'b0), .C(n14218), .Y(n14791) );
  NAND3X1 U2530 ( .A(n14398), .B(cs), .C(n34607), .Y(n14796) );
  OAI21X1 U2536 ( .A(n14802), .B(n14373), .C(n14803), .Y(n22522) );
  AOI21X1 U2537 ( .A(n30263), .B(1'b0), .C(n14218), .Y(n14803) );
  NAND3X1 U2541 ( .A(n14411), .B(cs), .C(n34607), .Y(n14808) );
  OAI21X1 U2547 ( .A(n14814), .B(n14373), .C(n14815), .Y(n22519) );
  AOI21X1 U2548 ( .A(n30258), .B(1'b0), .C(n14218), .Y(n14815) );
  NAND3X1 U2552 ( .A(n14424), .B(cs), .C(n34607), .Y(n14820) );
  OAI21X1 U2558 ( .A(n14826), .B(n14373), .C(n14827), .Y(n22516) );
  AOI21X1 U2559 ( .A(n30253), .B(1'b0), .C(n14218), .Y(n14827) );
  NAND3X1 U2563 ( .A(n14437), .B(cs), .C(n34607), .Y(n14832) );
  OAI21X1 U2569 ( .A(n14838), .B(n14373), .C(n14839), .Y(n22513) );
  AOI21X1 U2570 ( .A(n30248), .B(1'b0), .C(n14218), .Y(n14839) );
  NAND3X1 U2574 ( .A(n14450), .B(cs), .C(n34607), .Y(n14844) );
  OAI21X1 U2580 ( .A(n14850), .B(n14373), .C(n14851), .Y(n22510) );
  AOI21X1 U2581 ( .A(n30243), .B(1'b0), .C(n14218), .Y(n14851) );
  NAND3X1 U2585 ( .A(n14463), .B(cs), .C(n34607), .Y(n14856) );
  OAI21X1 U2591 ( .A(n14862), .B(n14373), .C(n14863), .Y(n22507) );
  AOI21X1 U2592 ( .A(n30238), .B(1'b0), .C(n14218), .Y(n14863) );
  NAND3X1 U2596 ( .A(n14476), .B(cs), .C(n34607), .Y(n14868) );
  NAND3X1 U2597 ( .A(n20812), .B(address[3]), .C(n24876), .Y(n14870) );
  OAI21X1 U2604 ( .A(n14876), .B(n14373), .C(n14877), .Y(n22504) );
  AOI21X1 U2605 ( .A(n30229), .B(1'b0), .C(n14218), .Y(n14877) );
  NAND3X1 U2609 ( .A(cs), .B(n14384), .C(n34605), .Y(n14882) );
  OAI21X1 U2615 ( .A(n14888), .B(n14373), .C(n14889), .Y(n22501) );
  AOI21X1 U2616 ( .A(n30220), .B(1'b0), .C(n14218), .Y(n14889) );
  NAND3X1 U2620 ( .A(n14398), .B(cs), .C(n34605), .Y(n14894) );
  OAI21X1 U2626 ( .A(n14900), .B(n14373), .C(n14901), .Y(n22498) );
  AOI21X1 U2627 ( .A(n30215), .B(1'b0), .C(n14218), .Y(n14901) );
  NAND3X1 U2631 ( .A(n14411), .B(cs), .C(n34605), .Y(n14906) );
  OAI21X1 U2637 ( .A(n14912), .B(n14373), .C(n14913), .Y(n22495) );
  AOI21X1 U2638 ( .A(n30210), .B(1'b0), .C(n14218), .Y(n14913) );
  NAND3X1 U2642 ( .A(n14424), .B(cs), .C(n34605), .Y(n14918) );
  OAI21X1 U2648 ( .A(n14924), .B(n14373), .C(n14925), .Y(n22492) );
  AOI21X1 U2649 ( .A(n30205), .B(1'b0), .C(n14218), .Y(n14925) );
  NAND3X1 U2653 ( .A(n14437), .B(cs), .C(n34605), .Y(n14930) );
  OAI21X1 U2659 ( .A(n14936), .B(n14373), .C(n14937), .Y(n22489) );
  AOI21X1 U2660 ( .A(n30200), .B(1'b0), .C(n14218), .Y(n14937) );
  NAND3X1 U2664 ( .A(n14450), .B(cs), .C(n34605), .Y(n14942) );
  OAI21X1 U2670 ( .A(n14948), .B(n14373), .C(n14949), .Y(n22486) );
  AOI21X1 U2671 ( .A(n30195), .B(1'b0), .C(n14218), .Y(n14949) );
  NAND3X1 U2675 ( .A(n14463), .B(cs), .C(n34605), .Y(n14954) );
  OAI21X1 U2681 ( .A(n14960), .B(n14373), .C(n14961), .Y(n22483) );
  AOI21X1 U2682 ( .A(n30190), .B(1'b0), .C(n14218), .Y(n14961) );
  NAND3X1 U2686 ( .A(n14476), .B(cs), .C(n34605), .Y(n14966) );
  NAND3X1 U2687 ( .A(n29469), .B(n34616), .C(n24875), .Y(n14968) );
  OAI21X1 U2694 ( .A(n14974), .B(n14373), .C(n14975), .Y(n22480) );
  AOI21X1 U2695 ( .A(n30180), .B(1'b0), .C(n14218), .Y(n14975) );
  NAND3X1 U2699 ( .A(cs), .B(n14384), .C(n34601), .Y(n14980) );
  OAI21X1 U2705 ( .A(n14986), .B(n14373), .C(n14987), .Y(n22477) );
  AOI21X1 U2706 ( .A(n30174), .B(1'b0), .C(n14218), .Y(n14987) );
  NAND3X1 U2710 ( .A(n14398), .B(cs), .C(n34601), .Y(n14992) );
  OAI21X1 U2716 ( .A(n14998), .B(n14373), .C(n14999), .Y(n22474) );
  AOI21X1 U2717 ( .A(n30169), .B(1'b0), .C(n14218), .Y(n14999) );
  NAND3X1 U2721 ( .A(n14411), .B(cs), .C(n34601), .Y(n15004) );
  OAI21X1 U2727 ( .A(n15010), .B(n14373), .C(n15011), .Y(n22471) );
  AOI21X1 U2728 ( .A(n30164), .B(1'b0), .C(n14218), .Y(n15011) );
  NAND3X1 U2732 ( .A(n14424), .B(cs), .C(n34601), .Y(n15016) );
  OAI21X1 U2738 ( .A(n15022), .B(n14373), .C(n15023), .Y(n22468) );
  AOI21X1 U2739 ( .A(n30159), .B(1'b0), .C(n14218), .Y(n15023) );
  NAND3X1 U2743 ( .A(n14437), .B(cs), .C(n34601), .Y(n15028) );
  OAI21X1 U2749 ( .A(n15034), .B(n14373), .C(n15035), .Y(n22465) );
  AOI21X1 U2750 ( .A(n30154), .B(1'b0), .C(n14218), .Y(n15035) );
  NAND3X1 U2754 ( .A(n14450), .B(cs), .C(n34601), .Y(n15040) );
  OAI21X1 U2760 ( .A(n15046), .B(n14373), .C(n15047), .Y(n22462) );
  AOI21X1 U2761 ( .A(n30149), .B(1'b0), .C(n14218), .Y(n15047) );
  NAND3X1 U2765 ( .A(n14463), .B(cs), .C(n34601), .Y(n15052) );
  OAI21X1 U2771 ( .A(n15058), .B(n14373), .C(n15059), .Y(n22459) );
  AOI21X1 U2772 ( .A(n30144), .B(1'b0), .C(n14218), .Y(n15059) );
  NAND3X1 U2776 ( .A(n14476), .B(cs), .C(n34601), .Y(n15064) );
  NAND3X1 U2777 ( .A(n34615), .B(n34616), .C(n26985), .Y(n15066) );
  OAI21X1 U2784 ( .A(n15071), .B(n14373), .C(n15072), .Y(n22456) );
  AOI21X1 U2785 ( .A(n30138), .B(1'b0), .C(n14218), .Y(n15072) );
  NAND3X1 U2789 ( .A(cs), .B(n14384), .C(n34598), .Y(n15077) );
  NOR3X1 U2790 ( .A(n29471), .B(n27715), .C(n29470), .Y(n14384) );
  OAI21X1 U2796 ( .A(n15083), .B(n14373), .C(n15084), .Y(n22453) );
  AOI21X1 U2797 ( .A(n30130), .B(1'b0), .C(n14218), .Y(n15084) );
  NAND3X1 U2801 ( .A(n14398), .B(cs), .C(n34598), .Y(n15089) );
  NOR3X1 U2802 ( .A(n29471), .B(n20978), .C(n29470), .Y(n14398) );
  OAI21X1 U2808 ( .A(n15095), .B(n14373), .C(n15096), .Y(n22450) );
  AOI21X1 U2809 ( .A(n30121), .B(1'b0), .C(n14218), .Y(n15096) );
  NAND3X1 U2813 ( .A(n14411), .B(cs), .C(n34598), .Y(n15101) );
  NOR3X1 U2814 ( .A(n27715), .B(n20811), .C(n29470), .Y(n14411) );
  OAI21X1 U2820 ( .A(n15107), .B(n14373), .C(n15108), .Y(n22447) );
  AOI21X1 U2821 ( .A(n30112), .B(1'b0), .C(n14218), .Y(n15108) );
  NAND3X1 U2825 ( .A(n14424), .B(cs), .C(n34598), .Y(n15113) );
  NOR3X1 U2826 ( .A(n20978), .B(n20811), .C(n29470), .Y(n14424) );
  OAI21X1 U2832 ( .A(n15119), .B(n14373), .C(n15120), .Y(n22444) );
  AOI21X1 U2833 ( .A(n30104), .B(1'b0), .C(n14218), .Y(n15120) );
  NAND3X1 U2837 ( .A(n14437), .B(cs), .C(n34598), .Y(n15125) );
  NOR3X1 U2838 ( .A(n27715), .B(n20810), .C(n29471), .Y(n14437) );
  OAI21X1 U2844 ( .A(n15131), .B(n14373), .C(n15132), .Y(n22441) );
  AOI21X1 U2845 ( .A(n30095), .B(1'b0), .C(n14218), .Y(n15132) );
  NAND3X1 U2849 ( .A(n14450), .B(cs), .C(n34598), .Y(n15137) );
  NOR3X1 U2850 ( .A(n20978), .B(n20810), .C(n29471), .Y(n14450) );
  OAI21X1 U2856 ( .A(n15143), .B(n14373), .C(n15144), .Y(n22438) );
  AOI21X1 U2857 ( .A(n30087), .B(1'b0), .C(n14218), .Y(n15144) );
  NAND3X1 U2861 ( .A(n14463), .B(cs), .C(n34598), .Y(n15149) );
  NOR3X1 U2862 ( .A(n20811), .B(n20810), .C(n27715), .Y(n14463) );
  OAI21X1 U2868 ( .A(n15156), .B(n14373), .C(n15157), .Y(n22435) );
  AOI21X1 U2869 ( .A(n30080), .B(1'b0), .C(n14218), .Y(n15157) );
  NAND3X1 U2874 ( .A(n14476), .B(cs), .C(n34598), .Y(n15167) );
  NAND3X1 U2875 ( .A(n34615), .B(n34616), .C(n27063), .Y(n15169) );
  NAND3X1 U2877 ( .A(n15170), .B(n15171), .C(n15172), .Y(n14675) );
  NOR3X1 U2878 ( .A(n24887), .B(n25108), .C(n24923), .Y(n15172) );
  NAND3X1 U2880 ( .A(data_in[6]), .B(n15177), .C(data_in[7]), .Y(n15173) );
  NOR3X1 U2881 ( .A(n15178), .B(n2264), .C(n2263), .Y(n15171) );
  NOR3X1 U2882 ( .A(address[7]), .B(n2262), .C(n2261), .Y(n15170) );
  NOR3X1 U2883 ( .A(n20811), .B(n20810), .C(n20978), .Y(n14476) );
  OAI21X1 U2885 ( .A(n25840), .B(n15180), .C(n15181), .Y(n22433) );
  OAI21X1 U2887 ( .A(n25760), .B(n15180), .C(n15185), .Y(n22432) );
  OAI21X1 U2889 ( .A(n25763), .B(n15180), .C(n15187), .Y(n22431) );
  OAI21X1 U2891 ( .A(n25663), .B(n15180), .C(n15189), .Y(n22430) );
  NAND3X1 U2895 ( .A(n23443), .B(n25210), .C(n15155), .Y(n15180) );
  AOI21X1 U2897 ( .A(n15155), .B(n24247), .C(n14218), .Y(n15195) );
  NAND2X1 U2901 ( .A(n15201), .B(n15202), .Y(n22428) );
  NAND3X1 U2902 ( .A(n34497), .B(n34614), .C(n34504), .Y(n15202) );
  OAI21X1 U2903 ( .A(n15204), .B(n22939), .C(n15201), .Y(n22427) );
  OAI21X1 U2904 ( .A(n15205), .B(n14373), .C(n15201), .Y(n22426) );
  OAI21X1 U2917 ( .A(n24277), .B(n14373), .C(n15201), .Y(n22425) );
  OAI21X1 U2930 ( .A(n15245), .B(n14373), .C(n15201), .Y(n22417) );
  NAND2X1 U2942 ( .A(n15201), .B(n15260), .Y(n22415) );
  OAI21X1 U2949 ( .A(n15269), .B(n14373), .C(n15201), .Y(n22414) );
  NAND2X1 U2962 ( .A(n15201), .B(n15283), .Y(n22412) );
  OAI21X1 U2969 ( .A(n15293), .B(n14373), .C(n15201), .Y(n22411) );
  NAND2X1 U2982 ( .A(n15201), .B(n15306), .Y(n22409) );
  OAI21X1 U2989 ( .A(n15316), .B(n14373), .C(n15201), .Y(n22408) );
  NAND2X1 U3002 ( .A(n15201), .B(n15329), .Y(n22406) );
  OAI21X1 U3009 ( .A(n15339), .B(n14373), .C(n15201), .Y(n22405) );
  NAND2X1 U3022 ( .A(n15201), .B(n15352), .Y(n22403) );
  OAI21X1 U3029 ( .A(n15362), .B(n14373), .C(n15201), .Y(n22402) );
  NAND2X1 U3042 ( .A(n15201), .B(n15377), .Y(n22400) );
  OAI21X1 U3049 ( .A(n15387), .B(n14373), .C(n15201), .Y(n22399) );
  NAND2X1 U3062 ( .A(n15201), .B(n15401), .Y(n22397) );
  OAI21X1 U3069 ( .A(n15411), .B(n14373), .C(n15201), .Y(n22396) );
  NAND2X1 U3082 ( .A(n15201), .B(n15424), .Y(n22394) );
  OAI21X1 U3089 ( .A(n15434), .B(n14373), .C(n15201), .Y(n22393) );
  NAND2X1 U3103 ( .A(n15201), .B(n15446), .Y(n22391) );
  OAI21X1 U3110 ( .A(n15456), .B(n14373), .C(n15201), .Y(n22390) );
  NAND2X1 U3124 ( .A(n15201), .B(n15469), .Y(n22388) );
  OAI21X1 U3131 ( .A(n15478), .B(n14373), .C(n15201), .Y(n22387) );
  NAND2X1 U3145 ( .A(n15201), .B(n15490), .Y(n22385) );
  OAI21X1 U3152 ( .A(n15500), .B(n14373), .C(n15201), .Y(n22384) );
  NAND2X1 U3166 ( .A(n15201), .B(n15512), .Y(n22382) );
  OAI21X1 U3173 ( .A(n15521), .B(n14373), .C(n15201), .Y(n22381) );
  OAI21X1 U3187 ( .A(n24275), .B(n14373), .C(n15201), .Y(n22379) );
  OAI21X1 U3194 ( .A(n15544), .B(n14373), .C(n15201), .Y(n22378) );
  OAI21X1 U3201 ( .A(n15552), .B(n14373), .C(n15201), .Y(n22377) );
  OAI21X1 U3212 ( .A(n24273), .B(n14373), .C(n15201), .Y(n22374) );
  NAND2X1 U3222 ( .A(n15201), .B(n15574), .Y(n22373) );
  OAI21X1 U3233 ( .A(n15589), .B(n14373), .C(n15201), .Y(n22371) );
  NAND2X1 U3246 ( .A(n15201), .B(n15601), .Y(n22369) );
  OAI21X1 U3254 ( .A(n15611), .B(n14373), .C(n15201), .Y(n22368) );
  NAND2X1 U3267 ( .A(n15201), .B(n15623), .Y(n22366) );
  OAI21X1 U3275 ( .A(n15632), .B(n14373), .C(n15201), .Y(n22365) );
  NAND2X1 U3288 ( .A(n15201), .B(n15644), .Y(n22363) );
  OAI21X1 U3296 ( .A(n15653), .B(n14373), .C(n15201), .Y(n22362) );
  NAND2X1 U3309 ( .A(n15201), .B(n15665), .Y(n22360) );
  OAI21X1 U3317 ( .A(n15674), .B(n14373), .C(n15201), .Y(n22359) );
  NAND2X1 U3330 ( .A(n15201), .B(n15686), .Y(n22357) );
  OAI21X1 U3338 ( .A(n15695), .B(n14373), .C(n15201), .Y(n22356) );
  NAND2X1 U3351 ( .A(n15201), .B(n15707), .Y(n22354) );
  OAI21X1 U3359 ( .A(n15716), .B(n14373), .C(n15201), .Y(n22353) );
  NAND2X1 U3372 ( .A(n15201), .B(n15729), .Y(n22351) );
  OAI21X1 U3380 ( .A(n15738), .B(n14373), .C(n15201), .Y(n22350) );
  NAND2X1 U3393 ( .A(n15201), .B(n15751), .Y(n22348) );
  OAI21X1 U3401 ( .A(n15760), .B(n14373), .C(n15201), .Y(n22347) );
  NAND2X1 U3414 ( .A(n15201), .B(n15772), .Y(n22345) );
  OAI21X1 U3422 ( .A(n15781), .B(n14373), .C(n15201), .Y(n22344) );
  NAND2X1 U3435 ( .A(n15201), .B(n15793), .Y(n22342) );
  OAI21X1 U3443 ( .A(n15802), .B(n14373), .C(n15201), .Y(n22341) );
  NAND2X1 U3456 ( .A(n15201), .B(n15814), .Y(n22339) );
  OAI21X1 U3464 ( .A(n15823), .B(n14373), .C(n15201), .Y(n22338) );
  NAND2X1 U3477 ( .A(n15201), .B(n15835), .Y(n22336) );
  OAI21X1 U3485 ( .A(n15844), .B(n14373), .C(n15201), .Y(n22335) );
  NAND2X1 U3498 ( .A(n15201), .B(n15856), .Y(n22333) );
  OAI21X1 U3506 ( .A(n15865), .B(n14373), .C(n15201), .Y(n22332) );
  NAND2X1 U3515 ( .A(n15201), .B(n15872), .Y(n22331) );
  NAND2X1 U3521 ( .A(n15201), .B(n15879), .Y(n22330) );
  OAI21X1 U3522 ( .A(n15873), .B(n15880), .C(n14097), .Y(n15879) );
  OAI21X1 U3529 ( .A(n15887), .B(n14373), .C(n15201), .Y(n22329) );
  OAI21X1 U3538 ( .A(n15897), .B(n14373), .C(n13994), .Y(n22328) );
  NAND2X1 U3540 ( .A(n15201), .B(n15899), .Y(n22327) );
  NAND2X1 U3541 ( .A(n14097), .B(n23904), .Y(n15899) );
  OAI21X1 U3551 ( .A(direct[0]), .B(n24692), .C(n15917), .Y(n15915) );
  OAI21X1 U3552 ( .A(n24278), .B(n24693), .C(direct[0]), .Y(n15917) );
  AOI21X1 U3554 ( .A(n15920), .B(n15921), .C(n24032), .Y(n15918) );
  AOI21X1 U3555 ( .A(n34568), .B(n15923), .C(n24031), .Y(n15922) );
  AOI21X1 U3556 ( .A(n34586), .B(n15925), .C(n24030), .Y(n15924) );
  AOI21X1 U3557 ( .A(n34589), .B(n15927), .C(n24020), .Y(n15926) );
  AOI22X1 U3558 ( .A(n15929), .B(n15930), .C(n34571), .D(n15931), .Y(n15928)
         );
  XNOR2X1 U3559 ( .A(n26917), .B(n25157), .Y(n15929) );
  FAX1 U3560 ( .A(n15934), .B(n15935), .C(n15936), .YC(), .YS(n15927) );
  FAX1 U3561 ( .A(n34569), .B(n15937), .C(n27185), .YC(), .YS(n15925) );
  FAX1 U3562 ( .A(n25146), .B(n27060), .C(n24987), .YC(), .YS(n15920) );
  AOI22X1 U3566 ( .A(n15937), .B(n15947), .C(n27185), .D(n34569), .Y(n15940)
         );
  AOI21X1 U3567 ( .A(n15935), .B(n15936), .C(n34570), .Y(n15938) );
  OAI21X1 U3568 ( .A(n15936), .B(n15935), .C(n15934), .Y(n15948) );
  OAI21X1 U3569 ( .A(n34576), .B(n15949), .C(n23896), .Y(n15934) );
  XNOR2X1 U3571 ( .A(n27096), .B(n27008), .Y(n15951) );
  XNOR2X1 U3572 ( .A(n27096), .B(n34574), .Y(n15949) );
  OAI21X1 U3575 ( .A(n25199), .B(n15956), .C(n23895), .Y(n15935) );
  XNOR2X1 U3577 ( .A(n27327), .B(n15955), .Y(n15958) );
  XNOR2X1 U3578 ( .A(n27327), .B(n26999), .Y(n15956) );
  OAI21X1 U3579 ( .A(n25199), .B(n15961), .C(n23887), .Y(n15960) );
  NAND3X1 U3580 ( .A(n15963), .B(n26930), .C(n24866), .Y(n15962) );
  AOI21X1 U3581 ( .A(n15955), .B(n26851), .C(n25200), .Y(n15965) );
  XNOR2X1 U3582 ( .A(n34573), .B(n34499), .Y(n15961) );
  NAND3X1 U3586 ( .A(n15970), .B(n26994), .C(n24865), .Y(n15943) );
  NAND3X1 U3587 ( .A(n27327), .B(n34499), .C(n15955), .Y(n15972) );
  NAND3X1 U3599 ( .A(n15979), .B(n26868), .C(n34575), .Y(n15978) );
  NAND3X1 U3600 ( .A(n15979), .B(n27177), .C(n24864), .Y(n15977) );
  AOI21X1 U3601 ( .A(n15953), .B(n26995), .C(n26868), .Y(n15982) );
  AOI21X1 U3602 ( .A(n24268), .B(n24255), .C(n34576), .Y(n15939) );
  NAND3X1 U3603 ( .A(n15987), .B(n26914), .C(n34577), .Y(n15980) );
  NOR3X1 U3604 ( .A(n27096), .B(n15979), .C(n27008), .Y(n15989) );
  AOI21X1 U3620 ( .A(n34506), .B(n34562), .C(n24029), .Y(n15916) );
  AOI21X1 U3621 ( .A(n15998), .B(n15921), .C(n24028), .Y(n15997) );
  AOI21X1 U3622 ( .A(n34563), .B(n15923), .C(n24027), .Y(n15999) );
  AOI21X1 U3623 ( .A(n34586), .B(n16001), .C(n26732), .Y(n16000) );
  AOI21X1 U3624 ( .A(n34589), .B(n16003), .C(n26733), .Y(n16002) );
  AOI22X1 U3625 ( .A(n16005), .B(n15930), .C(n34566), .D(n15931), .Y(n16004)
         );
  XNOR2X1 U3626 ( .A(n26918), .B(n26857), .Y(n16005) );
  FAX1 U3627 ( .A(n16008), .B(n16009), .C(n16010), .YC(), .YS(n16003) );
  FAX1 U3628 ( .A(n34564), .B(n16011), .C(n27006), .YC(), .YS(n16001) );
  FAX1 U3629 ( .A(n26854), .B(n26915), .C(n26749), .YC(), .YS(n15998) );
  AOI22X1 U3633 ( .A(n16011), .B(n16021), .C(n27006), .D(n34564), .Y(n16014)
         );
  AOI21X1 U3634 ( .A(n16009), .B(n16010), .C(n34565), .Y(n16012) );
  OAI21X1 U3635 ( .A(n16010), .B(n16009), .C(n16008), .Y(n16022) );
  OAI21X1 U3636 ( .A(n34596), .B(n16023), .C(n23894), .Y(n16008) );
  XNOR2X1 U3638 ( .A(n27182), .B(n27099), .Y(n16025) );
  XNOR2X1 U3639 ( .A(n27182), .B(n34594), .Y(n16023) );
  OAI21X1 U3642 ( .A(n34567), .B(n16030), .C(n26696), .Y(n16009) );
  XNOR2X1 U3644 ( .A(n27325), .B(n16187), .Y(n16032) );
  XNOR2X1 U3645 ( .A(n27325), .B(n27197), .Y(n16030) );
  OAI21X1 U3646 ( .A(n34567), .B(n16035), .C(n23886), .Y(n16034) );
  NAND3X1 U3647 ( .A(n16195), .B(n27193), .C(n24863), .Y(n16036) );
  AOI21X1 U3648 ( .A(n16187), .B(n27101), .C(n26859), .Y(n16039) );
  XNOR2X1 U3649 ( .A(n34501), .B(n34502), .Y(n16035) );
  NAND3X1 U3653 ( .A(n16044), .B(n27113), .C(n26920), .Y(n16017) );
  NAND3X1 U3666 ( .A(n16053), .B(n25219), .C(n34595), .Y(n16052) );
  NAND3X1 U3667 ( .A(n16053), .B(n27000), .C(n24862), .Y(n16051) );
  AOI21X1 U3668 ( .A(n16027), .B(n27076), .C(n25219), .Y(n16056) );
  AOI21X1 U3669 ( .A(n26855), .B(n26856), .C(n34596), .Y(n16013) );
  NOR3X1 U3671 ( .A(n27182), .B(n16053), .C(n27099), .Y(n16063) );
  AOI21X1 U3690 ( .A(n16075), .B(n15921), .C(n24026), .Y(n16073) );
  AOI21X1 U3691 ( .A(n34578), .B(n15923), .C(n24025), .Y(n16076) );
  AOI21X1 U3692 ( .A(n34586), .B(n16078), .C(n24024), .Y(n16077) );
  AOI21X1 U3693 ( .A(n34589), .B(n16080), .C(n24019), .Y(n16079) );
  AOI22X1 U3694 ( .A(n16082), .B(n15930), .C(n34581), .D(n15931), .Y(n16081)
         );
  XNOR2X1 U3695 ( .A(n25151), .B(n25156), .Y(n16082) );
  FAX1 U3696 ( .A(n16085), .B(n16086), .C(n16087), .YC(), .YS(n16080) );
  FAX1 U3697 ( .A(n34579), .B(n16088), .C(n27183), .YC(), .YS(n16078) );
  FAX1 U3698 ( .A(n25145), .B(n25119), .C(n24986), .YC(), .YS(n16075) );
  AOI22X1 U3702 ( .A(n16088), .B(n16098), .C(n27183), .D(n34579), .Y(n16091)
         );
  AOI21X1 U3703 ( .A(n16086), .B(n16087), .C(n34580), .Y(n16089) );
  OAI21X1 U3704 ( .A(n16087), .B(n16086), .C(n16085), .Y(n16099) );
  OAI21X1 U3705 ( .A(n23639), .B(n16100), .C(n23893), .Y(n16085) );
  XNOR2X1 U3707 ( .A(n27095), .B(n25422), .Y(n16102) );
  XNOR2X1 U3708 ( .A(n27095), .B(n34584), .Y(n16100) );
  OAI21X1 U3711 ( .A(n25197), .B(n16107), .C(n23892), .Y(n16086) );
  XNOR2X1 U3713 ( .A(n27326), .B(n16106), .Y(n16109) );
  XNOR2X1 U3714 ( .A(n27326), .B(n25341), .Y(n16107) );
  OAI21X1 U3715 ( .A(n25197), .B(n16112), .C(n23885), .Y(n16111) );
  NAND3X1 U3716 ( .A(n16114), .B(n27077), .C(n24861), .Y(n16113) );
  AOI21X1 U3717 ( .A(n16106), .B(n25113), .C(n25198), .Y(n16116) );
  XNOR2X1 U3718 ( .A(n34583), .B(n34500), .Y(n16112) );
  NAND3X1 U3722 ( .A(n16121), .B(n25207), .C(n24860), .Y(n16094) );
  NAND3X1 U3723 ( .A(n27326), .B(n34500), .C(n16106), .Y(n16123) );
  NAND3X1 U3735 ( .A(n16130), .B(n25216), .C(n34585), .Y(n16129) );
  NAND3X1 U3736 ( .A(n16130), .B(n26933), .C(n24859), .Y(n16128) );
  AOI21X1 U3737 ( .A(n16104), .B(n26867), .C(n25216), .Y(n16133) );
  AOI21X1 U3738 ( .A(n24267), .B(n24254), .C(n23639), .Y(n16090) );
  NOR3X1 U3740 ( .A(n27095), .B(n16130), .C(n25422), .Y(n16140) );
  AOI21X1 U3756 ( .A(n34506), .B(n34556), .C(n24023), .Y(n16071) );
  AOI21X1 U3757 ( .A(n16149), .B(n15921), .C(n24022), .Y(n16148) );
  AOI21X1 U3758 ( .A(n34557), .B(n15923), .C(n24021), .Y(n16150) );
  AOI21X1 U3759 ( .A(n34586), .B(n16152), .C(n26665), .Y(n16151) );
  AOI21X1 U3760 ( .A(n34589), .B(n16154), .C(n26666), .Y(n16153) );
  AOI22X1 U3761 ( .A(n16156), .B(n15930), .C(n34560), .D(n15931), .Y(n16155)
         );
  XOR2X1 U3762 ( .A(n26918), .B(n26858), .Y(n15930) );
  XNOR2X1 U3763 ( .A(n26918), .B(n26804), .Y(n16156) );
  FAX1 U3764 ( .A(n16161), .B(n16162), .C(n16163), .YC(), .YS(n16154) );
  FAX1 U3765 ( .A(n16164), .B(n16165), .C(n16166), .YC(), .YS(n15931) );
  FAX1 U3766 ( .A(n27085), .B(n27007), .C(n27184), .YC(), .YS(n15923) );
  FAX1 U3767 ( .A(n34558), .B(n16169), .C(n27097), .YC(), .YS(n16152) );
  FAX1 U3768 ( .A(n26801), .B(n26802), .C(n26800), .YC(), .YS(n16149) );
  AOI22X1 U3772 ( .A(n16169), .B(n16179), .C(n27097), .D(n34558), .Y(n16172)
         );
  AOI21X1 U3773 ( .A(n16162), .B(n16163), .C(n34559), .Y(n16170) );
  OAI21X1 U3774 ( .A(n16163), .B(n16162), .C(n16161), .Y(n16180) );
  OAI21X1 U3775 ( .A(n25214), .B(n16181), .C(n23891), .Y(n16161) );
  XNOR2X1 U3777 ( .A(n27005), .B(n27187), .Y(n16183) );
  XNOR2X1 U3778 ( .A(n27005), .B(n34591), .Y(n16181) );
  OAI21X1 U3781 ( .A(n34561), .B(n16188), .C(n26731), .Y(n16162) );
  XNOR2X1 U3783 ( .A(n27325), .B(n16187), .Y(n16190) );
  XNOR2X1 U3784 ( .A(n27325), .B(n27197), .Y(n16188) );
  OAI21X1 U3785 ( .A(n34561), .B(n16193), .C(n23884), .Y(n16192) );
  NAND3X1 U3786 ( .A(n16195), .B(n27193), .C(n24858), .Y(n16194) );
  AOI21X1 U3787 ( .A(n16187), .B(n27101), .C(n26919), .Y(n16197) );
  XNOR2X1 U3788 ( .A(n34501), .B(n34502), .Y(n16193) );
  NAND3X1 U3792 ( .A(n16202), .B(n27113), .C(n26920), .Y(n16175) );
  NAND3X1 U3793 ( .A(n27325), .B(n34502), .C(n16187), .Y(n16204) );
  NAND3X1 U3805 ( .A(n16211), .B(n25215), .C(n34592), .Y(n16210) );
  NAND3X1 U3806 ( .A(n16211), .B(n27086), .C(n24857), .Y(n16209) );
  AOI21X1 U3807 ( .A(n16185), .B(n26929), .C(n25215), .Y(n16214) );
  AOI21X1 U3808 ( .A(n26734), .B(n24253), .C(n25214), .Y(n16171) );
  NAND3X1 U3809 ( .A(n16219), .B(n26852), .C(n34593), .Y(n16212) );
  NOR3X1 U3810 ( .A(n27005), .B(n16211), .C(n27187), .Y(n16221) );
  XNOR2X1 U3826 ( .A(n26698), .B(n26699), .Y(n15921) );
  AOI22X1 U3827 ( .A(n27085), .B(n16231), .C(n27184), .D(n27007), .Y(n16230)
         );
  AOI21X1 U3828 ( .A(n16164), .B(n16166), .C(n34588), .Y(n16168) );
  OAI21X1 U3829 ( .A(n16166), .B(n16164), .C(n16165), .Y(n16232) );
  OAI21X1 U3830 ( .A(n16233), .B(n16234), .C(n26612), .Y(n16165) );
  OAI21X1 U3836 ( .A(n16242), .B(n16243), .C(n26638), .Y(n16164) );
  AOI21X1 U3840 ( .A(n16242), .B(n16247), .C(n34587), .Y(n16167) );
  OAI21X1 U3873 ( .A(n16269), .B(n14373), .C(n15201), .Y(n22325) );
  OAI21X1 U3882 ( .A(n16280), .B(n25080), .C(n15201), .Y(n22323) );
  NAND2X1 U3883 ( .A(reset), .B(n2219), .Y(n15201) );
  NAND2X1 U3885 ( .A(n14097), .B(n34505), .Y(n16280) );
  maze_router_DW01_add_9 r2497 ( .A(nc), .B({oc[31], n21116, oc[29:20], n26068, 
        oc[18:15], n25702, oc[13], n25709, oc[11:3], n21224, oc[1], n25692}), 
        .CI(1'b0), .SUM({n11685, n11684, n11683, n11682, n11681, n11680, 
        n11679, n11678, n11677, n11676, n11675, n11674, n11673, n11672, n11671, 
        n11670, n11669, n11668, n11667, n11666, n11665, n11664, n11663, n11662, 
        n11661, n11660, n11659, n11658, n11657, n11656, n11655, n11654}), 
        .CO() );
  maze_router_DW_mult_tc_2 r2498 ( .a(nc), .b({1'b0, 1'b1, 1'b1, 1'b0}), 
        .product({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, n11717, n11716, n11715, 
        n11714, n11713, n11712, n11711, n11710, n11709, n11708, n11707, n11706, 
        n11705, n11704, n11703, n11702, n11701, n11700, n11699, n11698, n11697, 
        n11696, n11695, n11694, n11693, n11692, n11691, n11690, n11689, n11688, 
        n11687, SYNOPSYS_UNCONNECTED_5}) );
  maze_router_DW01_add_10 r2500 ( .A({n11897, n11896, n11895, n11894, n11893, 
        n11892, n11891, n11890, n11889, n11888, n11887, n11886, n11885, n11884, 
        n11883, n11882, n11881, n11880, n11879, n11878, n11877, n11876, n11875, 
        n11874, n11873, n11872, n11871, n11870, n11869, n11868, n11867, n11866, 
        n11865, n11864, n11863, n11862, n11861, n11860, n11859, n11858, n11857, 
        n11856, n11855, n11854, n11853, n11852, n11851, n11850, n11849, n11848, 
        n11847, n11846, n11845, n11844, n11843, n11842, n11841, n11840, n11839, 
        n11838, n11837, n11836, n11835, n11834, n11833, n11832, n11831, n11830, 
        n11829, n11828, n11827, n11826, n11825, n11824, n11823, n11822, n11821, 
        n11820, n11819, n11818, n11817, n11816, n11815, n11814, n11813, n11812, 
        n11811, n11810, n11809, n11808, n11807, n11806, n11805, n11804, n11803, 
        n11802, n11801, n11800, n11799, n11798, n11797, n11796, n11795, n11794, 
        n11793, n11792, n11791, n11790, n11789, n11788, n11787, n11786, n11785, 
        n11784, n11783, n11782, n11781, n11780, n11779, n11778, n11777, n11776, 
        n11775, n11774, n11773, n11772, n11771, n11770, n11769, n11768, n11767, 
        n11766, n11765, n11764, n11763, n11762, n11761, n11760, n11759, n11758, 
        n11757, n11756, n11755, n11754, n11753, n11752, n11751, n11750, n11749, 
        n11748, n11747, n11746, n11745, n11744, n11743, n11742, n11741, n11740, 
        n11739, n11738, n11737, n11736, n11735, n11734, n11733, n11732, n11731, 
        n11730, n11729, n11728, n11727, n11726, n11725, n11724, n11723, n11722, 
        n11721, n11720, n11719, n11718}), .B({RN, n8229, n8228, n8227, n8226, 
        n8225, n8224, n8223, n8222, n8221, n8220, n8219, n8218, n8217, n8216, 
        n8215, n8214, n8213, n8212, n8211, n8210, n8209, n8208, n8207, n8206, 
        n8205, n8204, n8203, n8202, n8201, n8200, n8199, n8198, n8197, n8196, 
        n8195, n8194, n8193, n8192, n8191, n8190, n8189, n8188, n8187, n8186, 
        n8185, n8184, n8183, n8182, n8181, n8180, n8179, n8178, n8177, n8176, 
        n8175, n8174, n8173, n8172, n8171, n8170, n8169, n8168, n8167, n8166, 
        n8165, n8164, n8163, n8162, n8161, n8160, n8159, n8158, n8157, n8156, 
        n8155, n8154, n8153, n8152, n8151, n8150, n8149, n8148, n8147, n8146, 
        n8145, n8144, n8143, n8142, n8141, n8140, n8139, n8138, n8137, n8136, 
        n8135, n8134, n8133, n8132, n8131, n8130, n8129, n8128, n8127, n8126, 
        n8125, n8124, n8123, n8122, n8121, n8120, n8119, n8118, n8117, n8116, 
        n8115, n8114, n8113, n8112, n8111, n8110, n8109, n8108, n8107, n8106, 
        n8105, n8104, n8103, n8102, n8101, n8100, n8099, n8098, n8097, n8096, 
        n8095, n8094, n8093, n8092, n8091, n8090, n8089, n8088, n8087, n8086, 
        n8085, n8084, n8083, n8082, n8081, n8080, n8079, n8078, n8077, n8076, 
        n8075, n8074, n8073, n8072, n8071, n8070, n8069, n8068, n8067, n8066, 
        n8065, n8064, n8063, n8062, n8061, n8060, n8059, n8058, n8057, n8056}), 
        .CI(1'b0), .SUM({n12077, n12076, n12075, n12074, n12073, n12072, 
        n12071, n12070, n12069, n12068, n12067, n12066, n12065, n12064, n12063, 
        n12062, n12061, n12060, n12059, n12058, n12057, n12056, n12055, n12054, 
        n12053, n12052, n12051, n12050, n12049, n12048, n12047, n12046, n12045, 
        n12044, n12043, n12042, n12041, n12040, n12039, n12038, n12037, n12036, 
        n12035, n12034, n12033, n12032, n12031, n12030, n12029, n12028, n12027, 
        n12026, n12025, n12024, n12023, n12022, n12021, n12020, n12019, n12018, 
        n12017, n12016, n12015, n12014, n12013, n12012, n12011, n12010, n12009, 
        n12008, n12007, n12006, n12005, n12004, n12003, n12002, n12001, n12000, 
        n11999, n11998, n11997, n11996, n11995, n11994, n11993, n11992, n11991, 
        n11990, n11989, n11988, n11987, n11986, n11985, n11984, n11983, n11982, 
        n11981, n11980, n11979, n11978, n11977, n11976, n11975, n11974, n11973, 
        n11972, n11971, n11970, n11969, n11968, n11967, n11966, n11965, n11964, 
        n11963, n11962, n11961, n11960, n11959, n11958, n11957, n11956, n11955, 
        n11954, n11953, n11952, n11951, n11950, n11949, n11948, n11947, n11946, 
        n11945, n11944, n11943, n11942, n11941, n11940, n11939, n11938, n11937, 
        n11936, n11935, n11934, n11933, n11932, n11931, n11930, n11929, n11928, 
        n11927, n11926, n11925, n11924, n11923, n11922, n11921, n11920, n11919, 
        n11918, n11917, n11916, n11915, n11914, n11913, n11912, n11911, n11910, 
        n11909, n11908, n11907, n11906, n11905, n11904, n11903, n11902, n11901, 
        n11900, n11899, n11898}), .CO() );
  maze_router_DW01_dec_5 r2490 ( .A({oc[31], n21116, oc[29], n21140, n21141, 
        n26052, oc[25], n21118, oc[23], n21114, oc[21:20], n26068, n20968, 
        oc[17:15], n25702, oc[13], n25709, oc[11:3], n21224, oc[1], n25692}), 
        .SUM({n4221, n4220, n4219, n4218, n4217, n4216, n4215, n4214, n4213, 
        n4212, n4211, n4210, n4209, n4208, n4207, n4206, n4205, n4204, n4203, 
        n4202, n4201, n4200, n4199, n4198, n4197, n4196, n4195, n4194, n4193, 
        n4192, n4191, n4190}) );
  maze_router_DW01_inc_6 add_286 ( .A({nc[31:10], n25677, nc[8:7], n25612, 
        nc[5:4], n25718, n25613, nc[1:0]}), .SUM({n9157, n9156, n9155, n9154, 
        n9153, n9152, n9151, n9150, n9149, n9148, n9147, n9146, n9145, n9144, 
        n9143, n9142, n9141, n9140, n9139, n9138, n9137, n9136, n9135, n9134, 
        n9133, n9132, n9131, n9130, n9129, n9128, n9127, n9126}) );
  maze_router_DW01_inc_7 r2435 ( .A({oc[31], n21116, oc[29], n25573, n21141, 
        oc[26:23], n25646, oc[21:20], n26068, n20968, oc[17:15], n25713, 
        oc[13], n25709, oc[11:3], n21224, oc[1], n25692}), .SUM({n3307, n3306, 
        n3305, n3304, n3303, n3302, n3301, n3300, n3299, n3298, n3297, n3296, 
        n3295, n3294, n3293, n3292, n3291, n3290, n3289, n3288, n3287, n3286, 
        n3285, n3284, n3283, n3282, n3281, n3280, n3279, n3278, n3277, n3276})
         );
  maze_router_DW_leftsh_3 r2499 ( .A({RO, n3275, n3274, n3273, n3272, n3271, 
        n3270, n3269, n3268, n3267, n3266, n3265, n3264, n3263, n3262, n3261, 
        n3260, n3259, n3258, n3257, n3256, n3255, n3254, n3253, n3252, n3251, 
        n3250, n3249, n3248, n3247, n3246, n3245, n3244, n3243, n3242, n3241, 
        n3240, n3239, n3238, n3237, n3236, n3235, n3234, n3233, n3232, n3231, 
        n3230, n3229, n3228, n3227, n3226, n3225, n3224, n3223, n3222, n3221, 
        n3220, n3219, n3218, n3217, n3216, n3215, n3214, n3213, n3212, n3211, 
        n3210, n3209, n3208, n3207, n3206, n3205, n3204, n3203, n3202, n3201, 
        n3200, n3199, n3198, n3197, n3196, n3195, n3194, n3193, n3192, n3191, 
        n3190, n3189, n3188, n3187, n3186, n3185, n3184, n3183, n3182, n3181, 
        n3180, n3179, n3178, n3177, n3176, n3175, n3174, n3173, n3172, n3171, 
        n3170, n3169, n3168, n3167, n3166, n3165, n3164, n3163, n3162, n3161, 
        n3160, n3159, n3158, n3157, n3156, n3155, n3154, n3153, n3152, n3151, 
        n3150, n3149, n3148, n3147, n3146, n3145, n3144, n3143, n3142, n3141, 
        n3140, n3139, n3138, n3137, n3136, n3135, n3134, n3133, n3132, n3131, 
        n3130, n3129, n3128, n3127, n3126, n3125, n3124, n3123, n3122, n3121, 
        n3120, n3119, n3118, n3117, n3116, n3115, n3114, n3113, n3112, n3111, 
        n3110, n3109, n3108, n3107, n3106, n3105, n3104, n3103, n3102}), .SH({
        n11717, n11716, n11715, n11714, n11713, n11712, n11711, n11710, n11709, 
        n11708, n11707, n11706, n11705, n11704, n11703, n11702, n11701, n11700, 
        n11699, n11698, n11697, n11696, n11695, n11694, n11693, n11692, n11691, 
        n11690, n11689, n11688, n11687, 1'b0}), .B({n11897, n11896, n11895, 
        n11894, n11893, n11892, n11891, n11890, n11889, n11888, n11887, n11886, 
        n11885, n11884, n11883, n11882, n11881, n11880, n11879, n11878, n11877, 
        n11876, n11875, n11874, n11873, n11872, n11871, n11870, n11869, n11868, 
        n11867, n11866, n11865, n11864, n11863, n11862, n11861, n11860, n11859, 
        n11858, n11857, n11856, n11855, n11854, n11853, n11852, n11851, n11850, 
        n11849, n11848, n11847, n11846, n11845, n11844, n11843, n11842, n11841, 
        n11840, n11839, n11838, n11837, n11836, n11835, n11834, n11833, n11832, 
        n11831, n11830, n11829, n11828, n11827, n11826, n11825, n11824, n11823, 
        n11822, n11821, n11820, n11819, n11818, n11817, n11816, n11815, n11814, 
        n11813, n11812, n11811, n11810, n11809, n11808, n11807, n11806, n11805, 
        n11804, n11803, n11802, n11801, n11800, n11799, n11798, n11797, n11796, 
        n11795, n11794, n11793, n11792, n11791, n11790, n11789, n11788, n11787, 
        n11786, n11785, n11784, n11783, n11782, n11781, n11780, n11779, n11778, 
        n11777, n11776, n11775, n11774, n11773, n11772, n11771, n11770, n11769, 
        n11768, n11767, n11766, n11765, n11764, n11763, n11762, n11761, n11760, 
        n11759, n11758, n11757, n11756, n11755, n11754, n11753, n11752, n11751, 
        n11750, n11749, n11748, n11747, n11746, n11745, n11744, n11743, n11742, 
        n11741, n11740, n11739, n11738, n11737, n11736, n11735, n11734, n11733, 
        n11732, n11731, n11730, n11729, n11728, n11727, n11726, n11725, n11724, 
        n11723, n11722, n11721, n11720, n11719, n11718}) );
  AND2X2 U8518 ( .A(n23285), .B(n32491), .Y(n20806) );
  INVX1 U8519 ( .A(net151801), .Y(n20807) );
  BUFX2 U8520 ( .A(n26049), .Y(n20808) );
  INVX1 U8521 ( .A(n29463), .Y(n20809) );
  INVX1 U8522 ( .A(n29470), .Y(n20810) );
  INVX4 U8523 ( .A(n8052), .Y(n29463) );
  INVX1 U8524 ( .A(n29471), .Y(n20811) );
  BUFX2 U8525 ( .A(address[4]), .Y(n20812) );
  INVX1 U8526 ( .A(n2256), .Y(n29508) );
  OR2X2 U8527 ( .A(n29580), .B(n21168), .Y(n29581) );
  INVX1 U8528 ( .A(alt5_net95670), .Y(n20813) );
  INVX4 U8529 ( .A(n2251), .Y(alt5_net95670) );
  INVX1 U8530 ( .A(alt5_net95668), .Y(n20872) );
  AND2X2 U8531 ( .A(net90053), .B(n20814), .Y(n32197) );
  AND2X2 U8532 ( .A(n29704), .B(net96340), .Y(n20814) );
  INVX4 U8533 ( .A(n30078), .Y(n29353) );
  MUX2X1 U8534 ( .B(n29166), .A(n29165), .S(n29179), .Y(n29164) );
  INVX4 U8535 ( .A(n29179), .Y(n29180) );
  INVX1 U8536 ( .A(n31921), .Y(n20815) );
  INVX1 U8537 ( .A(n31921), .Y(n20816) );
  INVX1 U8538 ( .A(n31921), .Y(n20817) );
  INVX1 U8539 ( .A(n31921), .Y(n32099) );
  INVX1 U8540 ( .A(n26056), .Y(n20818) );
  INVX1 U8541 ( .A(n29209), .Y(n20819) );
  INVX1 U8542 ( .A(n29209), .Y(n20820) );
  INVX4 U8543 ( .A(n29209), .Y(n29235) );
  BUFX2 U8544 ( .A(n26448), .Y(n20821) );
  INVX1 U8545 ( .A(n29314), .Y(n20822) );
  INVX1 U8546 ( .A(n27299), .Y(n29231) );
  INVX1 U8547 ( .A(n31921), .Y(n20823) );
  INVX1 U8548 ( .A(n29236), .Y(n20824) );
  INVX1 U8549 ( .A(n29236), .Y(n20825) );
  INVX1 U8550 ( .A(n29236), .Y(n29234) );
  INVX2 U8551 ( .A(n27299), .Y(n26463) );
  INVX2 U8552 ( .A(n27299), .Y(n26464) );
  INVX4 U8553 ( .A(n29253), .Y(n26310) );
  INVX1 U8554 ( .A(n29236), .Y(n20826) );
  INVX1 U8555 ( .A(n29236), .Y(n20827) );
  INVX1 U8556 ( .A(n25184), .Y(n20828) );
  INVX2 U8557 ( .A(n30707), .Y(n25184) );
  INVX1 U8558 ( .A(n29236), .Y(n20829) );
  BUFX2 U8559 ( .A(n31901), .Y(n29208) );
  INVX2 U8560 ( .A(n29204), .Y(n29236) );
  INVX2 U8561 ( .A(n30928), .Y(n23011) );
  OR2X1 U8562 ( .A(n31661), .B(n31668), .Y(n31669) );
  INVX1 U8563 ( .A(n30727), .Y(n25185) );
  AND2X1 U8564 ( .A(n30716), .B(net96340), .Y(n30727) );
  OR2X2 U8565 ( .A(n23245), .B(n31095), .Y(n20830) );
  BUFX2 U8566 ( .A(grid[223]), .Y(n20831) );
  OR2X2 U8567 ( .A(n23221), .B(n20832), .Y(n23220) );
  OR2X1 U8568 ( .A(n30738), .B(n23222), .Y(n20832) );
  INVX1 U8569 ( .A(n23081), .Y(n20833) );
  AND2X1 U8570 ( .A(n31444), .B(net96340), .Y(n31454) );
  INVX1 U8571 ( .A(n26278), .Y(n20834) );
  OR2X2 U8572 ( .A(n23619), .B(n30939), .Y(n20835) );
  INVX2 U8573 ( .A(n31334), .Y(n23036) );
  INVX2 U8574 ( .A(n31803), .Y(n23061) );
  OAI21X1 U8575 ( .A(n20837), .B(net96592), .C(n20838), .Y(n20836) );
  INVX1 U8576 ( .A(n20836), .Y(n33521) );
  INVX8 U8577 ( .A(n12002), .Y(n20837) );
  INVX8 U8578 ( .A(n33519), .Y(n20838) );
  INVX4 U8579 ( .A(net96592), .Y(net96574) );
  INVX1 U8580 ( .A(n26278), .Y(n20839) );
  INVX1 U8581 ( .A(n26278), .Y(n20840) );
  INVX1 U8582 ( .A(n31162), .Y(n20841) );
  MUX2X1 U8583 ( .B(n28687), .A(n28690), .S(n20842), .Y(n28701) );
  INVX8 U8584 ( .A(n26555), .Y(n20842) );
  INVX1 U8585 ( .A(n26294), .Y(n20843) );
  INVX1 U8586 ( .A(n31280), .Y(n20844) );
  BUFX2 U8587 ( .A(grid[301]), .Y(n20845) );
  INVX2 U8588 ( .A(n26292), .Y(n26294) );
  AND2X2 U8589 ( .A(n21529), .B(n24881), .Y(n32641) );
  INVX2 U8590 ( .A(n26517), .Y(n26146) );
  AND2X2 U8591 ( .A(n27159), .B(n25458), .Y(n21176) );
  MUX2X1 U8592 ( .B(n28584), .A(n28585), .S(n20846), .Y(n28583) );
  INVX8 U8593 ( .A(n21075), .Y(n20846) );
  INVX1 U8594 ( .A(n21097), .Y(n20847) );
  INVX1 U8595 ( .A(n25079), .Y(n20848) );
  INVX1 U8596 ( .A(n28598), .Y(n20849) );
  INVX2 U8597 ( .A(n27904), .Y(n20850) );
  INVX4 U8598 ( .A(n25679), .Y(n27910) );
  INVX2 U8599 ( .A(n25860), .Y(n34406) );
  INVX4 U8600 ( .A(net96604), .Y(net96576) );
  INVX1 U8601 ( .A(net107076), .Y(n20851) );
  XNOR2X1 U8602 ( .A(n34238), .B(n20852), .Y(n26057) );
  INVX8 U8603 ( .A(n34239), .Y(n20852) );
  INVX1 U8604 ( .A(net116755), .Y(n20853) );
  INVX4 U8605 ( .A(n33661), .Y(n27207) );
  INVX4 U8606 ( .A(n33215), .Y(n21387) );
  INVX4 U8607 ( .A(n33398), .Y(n21384) );
  INVX2 U8608 ( .A(n33276), .Y(n25430) );
  INVX4 U8609 ( .A(n33470), .Y(n25427) );
  INVX2 U8610 ( .A(n33726), .Y(n26764) );
  INVX8 U8611 ( .A(n23111), .Y(n33762) );
  INVX4 U8612 ( .A(n33747), .Y(n23111) );
  INVX4 U8613 ( .A(n33770), .Y(n21378) );
  INVX4 U8614 ( .A(n33837), .Y(n21375) );
  INVX2 U8615 ( .A(n22970), .Y(n23467) );
  INVX8 U8616 ( .A(n23110), .Y(n33884) );
  INVX4 U8617 ( .A(n29760), .Y(n23110) );
  INVX4 U8618 ( .A(n25203), .Y(n33538) );
  INVX4 U8619 ( .A(n32910), .Y(n25452) );
  INVX4 U8620 ( .A(n29190), .Y(n32773) );
  INVX8 U8621 ( .A(n25347), .Y(n33471) );
  INVX2 U8622 ( .A(n21174), .Y(n25347) );
  INVX4 U8623 ( .A(n32895), .Y(n26269) );
  INVX2 U8624 ( .A(n32913), .Y(n25454) );
  INVX8 U8625 ( .A(n23112), .Y(n33247) );
  INVX4 U8626 ( .A(n32518), .Y(n23112) );
  INVX4 U8627 ( .A(n29373), .Y(n29371) );
  INVX8 U8628 ( .A(n29372), .Y(n29370) );
  INVX2 U8629 ( .A(n21162), .Y(n29385) );
  INVX2 U8630 ( .A(net96586), .Y(net96558) );
  INVX4 U8631 ( .A(net96600), .Y(net96588) );
  INVX4 U8632 ( .A(net102091), .Y(net96604) );
  INVX2 U8633 ( .A(net96598), .Y(net96584) );
  INVX2 U8634 ( .A(n26325), .Y(n26327) );
  INVX2 U8635 ( .A(n31883), .Y(n23210) );
  INVX2 U8636 ( .A(n31661), .Y(n23050) );
  AND2X2 U8637 ( .A(net96340), .B(n31654), .Y(n31661) );
  INVX2 U8638 ( .A(n31274), .Y(n23033) );
  AND2X2 U8639 ( .A(n31267), .B(net96340), .Y(n31274) );
  INVX2 U8640 ( .A(n34442), .Y(n25619) );
  INVX4 U8641 ( .A(n25619), .Y(n34355) );
  INVX2 U8642 ( .A(n25661), .Y(n27912) );
  INVX2 U8643 ( .A(n34443), .Y(n25620) );
  INVX2 U8644 ( .A(n33111), .Y(n23093) );
  INVX4 U8645 ( .A(n34309), .Y(n34323) );
  INVX4 U8646 ( .A(n23427), .Y(n25446) );
  AND2X2 U8647 ( .A(n34291), .B(n34351), .Y(n34311) );
  INVX4 U8648 ( .A(n22962), .Y(n33158) );
  AND2X2 U8649 ( .A(n34322), .B(n34309), .Y(n34320) );
  AND2X2 U8650 ( .A(n31868), .B(n23443), .Y(n27261) );
  INVX2 U8651 ( .A(n29270), .Y(n29268) );
  AND2X2 U8652 ( .A(n31868), .B(n27304), .Y(n27271) );
  INVX2 U8653 ( .A(n27262), .Y(n29312) );
  INVX4 U8654 ( .A(n29347), .Y(n29343) );
  INVX4 U8655 ( .A(n29343), .Y(n29351) );
  INVX4 U8656 ( .A(n29443), .Y(n28220) );
  INVX1 U8657 ( .A(net53596), .Y(net149982) );
  INVX2 U8658 ( .A(n29357), .Y(n29355) );
  INVX2 U8659 ( .A(alt14_net96326), .Y(net105813) );
  INVX2 U8660 ( .A(alt14_net96328), .Y(net105814) );
  INVX2 U8661 ( .A(alt14_net96326), .Y(net105810) );
  INVX8 U8662 ( .A(net104479), .Y(net53601) );
  INVX8 U8663 ( .A(net89785), .Y(net104479) );
  INVX1 U8664 ( .A(n25163), .Y(n32266) );
  INVX2 U8665 ( .A(n29253), .Y(n26314) );
  INVX2 U8666 ( .A(n29253), .Y(n26307) );
  INVX4 U8667 ( .A(n27276), .Y(n29253) );
  INVX2 U8668 ( .A(n25782), .Y(n25821) );
  INVX1 U8669 ( .A(net151812), .Y(n20854) );
  INVX1 U8670 ( .A(net109766), .Y(n20855) );
  INVX2 U8671 ( .A(net113687), .Y(net105803) );
  MUX2X1 U8672 ( .B(grid[185]), .A(grid[191]), .S(net150251), .Y(n20905) );
  MUX2X1 U8673 ( .B(n28060), .A(n28059), .S(net147761), .Y(n28058) );
  INVX1 U8674 ( .A(n34290), .Y(n34291) );
  INVX4 U8675 ( .A(n21131), .Y(n34305) );
  AND2X2 U8676 ( .A(n32996), .B(n32995), .Y(n32997) );
  INVX1 U8677 ( .A(n25349), .Y(n20856) );
  INVX2 U8678 ( .A(n34262), .Y(n25689) );
  INVX4 U8679 ( .A(n25349), .Y(n33912) );
  XNOR2X1 U8680 ( .A(n21113), .B(n20857), .Y(n34270) );
  XNOR2X1 U8681 ( .A(n25759), .B(n34264), .Y(n20857) );
  AND2X2 U8682 ( .A(n3270), .B(n33216), .Y(n20858) );
  AND2X2 U8683 ( .A(n3264), .B(n33247), .Y(n20859) );
  NOR2X1 U8684 ( .A(n20858), .B(n20859), .Y(n32707) );
  INVX1 U8685 ( .A(n20964), .Y(n34329) );
  INVX1 U8686 ( .A(net143105), .Y(n4126) );
  BUFX2 U8687 ( .A(net95482), .Y(net143105) );
  INVX1 U8688 ( .A(n4126), .Y(net108471) );
  INVX1 U8689 ( .A(n4126), .Y(net95477) );
  AOI21X1 U8690 ( .A(direction_line[1]), .B(n20865), .C(net145121), .Y(
        net95482) );
  INVX1 U8691 ( .A(n20863), .Y(n20865) );
  OR2X2 U8692 ( .A(n20864), .B(net143109), .Y(n20863) );
  INVX1 U8693 ( .A(net53176), .Y(net145121) );
  INVX1 U8694 ( .A(net143105), .Y(net115619) );
  OR2X2 U8695 ( .A(n20866), .B(n20867), .Y(n20864) );
  OR2X2 U8696 ( .A(net110927), .B(net114253), .Y(n20866) );
  INVX1 U8697 ( .A(net110926), .Y(net110927) );
  INVX1 U8698 ( .A(net114252), .Y(net114253) );
  AND2X2 U8699 ( .A(n20860), .B(pLoc[1]), .Y(n20867) );
  AND2X2 U8700 ( .A(n20861), .B(n20862), .Y(n20860) );
  INVX1 U8701 ( .A(net111628), .Y(net143109) );
  INVX1 U8702 ( .A(n20863), .Y(net145295) );
  INVX1 U8703 ( .A(pLoc[2]), .Y(n20861) );
  INVX1 U8704 ( .A(pLoc[3]), .Y(n20862) );
  AND2X2 U8705 ( .A(n20860), .B(pLoc[1]), .Y(net109417) );
  INVX8 U8706 ( .A(alt14_net96276), .Y(alt14_net96264) );
  INVX4 U8707 ( .A(net105988), .Y(alt14_net96276) );
  INVX1 U8708 ( .A(net90064), .Y(net105988) );
  INVX1 U8709 ( .A(alt14_net96276), .Y(net112192) );
  INVX1 U8710 ( .A(alt14_net96276), .Y(net111237) );
  INVX4 U8711 ( .A(alt14_net96276), .Y(net109766) );
  MUX2X1 U8712 ( .B(n20869), .A(net111984), .S(n20872), .Y(net90064) );
  AND2X2 U8713 ( .A(net143040), .B(n20871), .Y(n20869) );
  BUFX2 U8714 ( .A(n14360), .Y(net143040) );
  BUFX2 U8715 ( .A(n14359), .Y(n20871) );
  NAND3X1 U8716 ( .A(n20868), .B(net111332), .C(net139028), .Y(n14359) );
  INVX1 U8717 ( .A(net149764), .Y(n20868) );
  AND2X2 U8718 ( .A(net146826), .B(net109440), .Y(net149764) );
  AND2X2 U8719 ( .A(net142789), .B(net109485), .Y(net111332) );
  INVX1 U8720 ( .A(net108471), .Y(net139028) );
  AND2X2 U8721 ( .A(net114808), .B(net143010), .Y(net111984) );
  INVX4 U8722 ( .A(n2251), .Y(alt5_net95668) );
  INVX1 U8723 ( .A(net105988), .Y(alt14_net96258) );
  NAND3X1 U8724 ( .A(net109385), .B(n20870), .C(net95477), .Y(n14360) );
  AND2X2 U8725 ( .A(net109440), .B(net146826), .Y(net109385) );
  INVX1 U8726 ( .A(net108478), .Y(n20870) );
  AND2X2 U8727 ( .A(net142788), .B(net109485), .Y(net108478) );
  INVX1 U8728 ( .A(net143040), .Y(net94649) );
  BUFX2 U8729 ( .A(net90056), .Y(net142746) );
  NAND3X1 U8730 ( .A(net108803), .B(net110685), .C(n20939), .Y(net90056) );
  MUX2X1 U8731 ( .B(net108805), .A(net108804), .S(net110421), .Y(net108803) );
  MUX2X1 U8732 ( .B(net110687), .A(net110686), .S(net110421), .Y(net110685) );
  NOR3X1 U8733 ( .A(net114723), .B(n20940), .C(n20938), .Y(n20939) );
  INVX1 U8734 ( .A(n4227), .Y(net114723) );
  INVX1 U8735 ( .A(n4226), .Y(n20940) );
  MUX2X1 U8736 ( .B(alt14_net6129), .A(alt14_net6130), .S(net110421), .Y(n4226) );
  AND2X2 U8737 ( .A(n20941), .B(n4223), .Y(n20938) );
  INVX1 U8738 ( .A(net142746), .Y(net147735) );
  INVX1 U8739 ( .A(net142746), .Y(net151709) );
  INVX1 U8740 ( .A(n4224), .Y(n20941) );
  MUX2X1 U8741 ( .B(alt14_net6254), .A(alt14_net6253), .S(net53623), .Y(n4224)
         );
  MUX2X1 U8742 ( .B(n20934), .A(n20933), .S(net53623), .Y(n4223) );
  BUFX2 U8743 ( .A(n20938), .Y(net108311) );
  MUX2X1 U8744 ( .B(n20885), .A(n20900), .S(net89785), .Y(n20934) );
  MUX2X1 U8745 ( .B(n20886), .A(n20887), .S(net113954), .Y(n20885) );
  MUX2X1 U8746 ( .B(n20882), .A(n20879), .S(net150245), .Y(n20886) );
  MUX2X1 U8747 ( .B(n20884), .A(n20883), .S(net105821), .Y(n20882) );
  MUX2X1 U8748 ( .B(grid[305]), .A(grid[311]), .S(alt14_net96248), .Y(n20884)
         );
  INVX1 U8749 ( .A(alt14_net96268), .Y(alt14_net96248) );
  MUX2X1 U8750 ( .B(grid[293]), .A(grid[299]), .S(alt14_net96248), .Y(n20883)
         );
  INVX2 U8751 ( .A(net113686), .Y(net105821) );
  MUX2X1 U8752 ( .B(n20880), .A(n20881), .S(net105795), .Y(n20879) );
  MUX2X1 U8753 ( .B(grid[317]), .A(grid[323]), .S(net111205), .Y(n20880) );
  INVX1 U8754 ( .A(alt14_net96268), .Y(net111205) );
  MUX2X1 U8755 ( .B(grid[329]), .A(grid[335]), .S(net105787), .Y(n20881) );
  INVX8 U8756 ( .A(alt14_net96264), .Y(net105787) );
  INVX1 U8757 ( .A(net115636), .Y(net105795) );
  INVX1 U8758 ( .A(alt14_net96302), .Y(net150245) );
  MUX2X1 U8759 ( .B(n20876), .A(n20873), .S(net149982), .Y(n20887) );
  MUX2X1 U8760 ( .B(n20877), .A(n20878), .S(net105796), .Y(n20876) );
  MUX2X1 U8761 ( .B(grid[341]), .A(grid[347]), .S(alt14_net96230), .Y(n20877)
         );
  INVX8 U8762 ( .A(alt14_net96264), .Y(alt14_net96230) );
  MUX2X1 U8763 ( .B(grid[353]), .A(grid[359]), .S(net112202), .Y(n20878) );
  INVX8 U8764 ( .A(net105786), .Y(net112202) );
  INVX1 U8765 ( .A(net115636), .Y(net105796) );
  MUX2X1 U8766 ( .B(n20874), .A(n20875), .S(net105810), .Y(n20873) );
  MUX2X1 U8767 ( .B(grid[365]), .A(grid[371]), .S(alt14_net96230), .Y(n20874)
         );
  MUX2X1 U8768 ( .B(grid[377]), .A(grid[383]), .S(alt14_net96236), .Y(n20875)
         );
  INVX8 U8769 ( .A(alt14_net96264), .Y(alt14_net96236) );
  OAI21X1 U8770 ( .A(net110410), .B(net89744), .C(net142478), .Y(net113954) );
  MUX2X1 U8771 ( .B(n20901), .A(n20902), .S(net113955), .Y(n20900) );
  MUX2X1 U8772 ( .B(n20897), .A(n20894), .S(n20935), .Y(n20901) );
  MUX2X1 U8773 ( .B(n20898), .A(n20899), .S(net105810), .Y(n20897) );
  MUX2X1 U8774 ( .B(grid[203]), .A(grid[197]), .S(net109766), .Y(n20898) );
  MUX2X1 U8775 ( .B(grid[209]), .A(grid[215]), .S(net105787), .Y(n20899) );
  MUX2X1 U8776 ( .B(n20895), .A(n20896), .S(net105799), .Y(n20894) );
  MUX2X1 U8777 ( .B(grid[221]), .A(grid[227]), .S(net111205), .Y(n20895) );
  INVX1 U8778 ( .A(net111237), .Y(net149909) );
  MUX2X1 U8779 ( .B(grid[233]), .A(grid[239]), .S(net105787), .Y(n20896) );
  INVX1 U8780 ( .A(net115636), .Y(net105799) );
  INVX1 U8781 ( .A(alt14_net96304), .Y(n20935) );
  MUX2X1 U8782 ( .B(n20891), .A(n20888), .S(net149936), .Y(n20902) );
  MUX2X1 U8783 ( .B(n20892), .A(n20893), .S(net105814), .Y(n20891) );
  MUX2X1 U8784 ( .B(grid[245]), .A(grid[251]), .S(net150261), .Y(n20892) );
  INVX1 U8785 ( .A(alt14_net96264), .Y(net150261) );
  MUX2X1 U8786 ( .B(grid[263]), .A(grid[257]), .S(net137490), .Y(n20893) );
  INVX4 U8787 ( .A(net137489), .Y(net137490) );
  MUX2X1 U8788 ( .B(n20889), .A(n20890), .S(net105813), .Y(n20888) );
  MUX2X1 U8789 ( .B(grid[269]), .A(grid[275]), .S(net105787), .Y(n20889) );
  MUX2X1 U8790 ( .B(grid[287]), .A(grid[281]), .S(net115535), .Y(n20890) );
  INVX1 U8791 ( .A(net112188), .Y(net115535) );
  INVX8 U8792 ( .A(net53596), .Y(net149936) );
  OAI21X1 U8793 ( .A(net110410), .B(net89744), .C(net142478), .Y(net113955) );
  AND2X2 U8794 ( .A(net104480), .B(net95457), .Y(net89785) );
  MUX2X1 U8795 ( .B(n20930), .A(n20915), .S(net104479), .Y(n20933) );
  MUX2X1 U8796 ( .B(n20931), .A(n20932), .S(net113954), .Y(n20930) );
  MUX2X1 U8797 ( .B(n20927), .A(n20924), .S(net149986), .Y(n20931) );
  MUX2X1 U8798 ( .B(n20929), .A(n20928), .S(net149877), .Y(n20927) );
  MUX2X1 U8799 ( .B(grid[17]), .A(grid[23]), .S(alt14_net96230), .Y(n20929) );
  MUX2X1 U8800 ( .B(grid[5]), .A(grid[11]), .S(alt14_net96236), .Y(n20928) );
  INVX1 U8801 ( .A(net115635), .Y(net149877) );
  MUX2X1 U8802 ( .B(n20925), .A(n20926), .S(net105813), .Y(n20924) );
  MUX2X1 U8803 ( .B(grid[29]), .A(grid[35]), .S(net150261), .Y(n20925) );
  MUX2X1 U8804 ( .B(grid[47]), .A(grid[41]), .S(net137490), .Y(n20926) );
  INVX2 U8805 ( .A(alt14_net96304), .Y(net149986) );
  MUX2X1 U8806 ( .B(n20918), .A(n20921), .S(n20936), .Y(n20932) );
  MUX2X1 U8807 ( .B(n20919), .A(n20920), .S(net105815), .Y(n20918) );
  MUX2X1 U8808 ( .B(grid[77]), .A(grid[83]), .S(alt14_net96236), .Y(n20919) );
  MUX2X1 U8809 ( .B(grid[95]), .A(grid[89]), .S(net105778), .Y(n20920) );
  INVX4 U8810 ( .A(alt14_net96250), .Y(net105778) );
  INVX1 U8811 ( .A(net149876), .Y(net105815) );
  MUX2X1 U8812 ( .B(n20923), .A(n20922), .S(net113687), .Y(n20921) );
  MUX2X1 U8813 ( .B(grid[65]), .A(grid[71]), .S(net112202), .Y(n20923) );
  MUX2X1 U8814 ( .B(grid[53]), .A(grid[59]), .S(net110246), .Y(n20922) );
  INVX4 U8815 ( .A(net105786), .Y(net110246) );
  INVX4 U8816 ( .A(net113686), .Y(net113687) );
  INVX1 U8817 ( .A(net150245), .Y(n20936) );
  MUX2X1 U8818 ( .B(n20917), .A(n20916), .S(n20937), .Y(n20915) );
  MUX2X1 U8819 ( .B(n20906), .A(n20903), .S(net149986), .Y(n20917) );
  MUX2X1 U8820 ( .B(n20907), .A(n20908), .S(net105810), .Y(n20906) );
  MUX2X1 U8821 ( .B(grid[149]), .A(grid[155]), .S(net105787), .Y(n20907) );
  MUX2X1 U8822 ( .B(grid[161]), .A(grid[167]), .S(net112202), .Y(n20908) );
  MUX2X1 U8823 ( .B(n20904), .A(n20905), .S(net105814), .Y(n20903) );
  MUX2X1 U8824 ( .B(grid[173]), .A(grid[179]), .S(n20855), .Y(n20904) );
  INVX1 U8825 ( .A(net112188), .Y(net116755) );
  MUX2X1 U8826 ( .B(n20909), .A(n20912), .S(net114744), .Y(n20916) );
  MUX2X1 U8827 ( .B(n20910), .A(n20911), .S(net105807), .Y(n20909) );
  MUX2X1 U8828 ( .B(grid[125]), .A(grid[131]), .S(net112202), .Y(n20910) );
  MUX2X1 U8829 ( .B(grid[137]), .A(grid[143]), .S(n20853), .Y(n20911) );
  INVX1 U8830 ( .A(alt14_net96326), .Y(net105807) );
  MUX2X1 U8831 ( .B(n20913), .A(n20914), .S(net105798), .Y(n20912) );
  MUX2X1 U8832 ( .B(grid[101]), .A(grid[107]), .S(net112202), .Y(n20913) );
  MUX2X1 U8833 ( .B(grid[113]), .A(grid[119]), .S(alt14_net96236), .Y(n20914)
         );
  INVX4 U8834 ( .A(net113687), .Y(net105798) );
  INVX1 U8835 ( .A(n20935), .Y(net114744) );
  INVX1 U8836 ( .A(net113955), .Y(n20937) );
  INVX4 U8837 ( .A(net124029), .Y(net53623) );
  BUFX2 U8838 ( .A(n4223), .Y(net149850) );
  INVX1 U8839 ( .A(n21834), .Y(net146640) );
  AND2X2 U8840 ( .A(n20945), .B(n20947), .Y(n21834) );
  INVX1 U8841 ( .A(n20949), .Y(n20945) );
  AND2X2 U8842 ( .A(n11672), .B(net96576), .Y(n20949) );
  BUFX2 U8843 ( .A(n20948), .Y(n20947) );
  AOI22X1 U8844 ( .A(n4208), .B(net147506), .C(n3294), .D(n20942), .Y(n20948)
         );
  INVX1 U8845 ( .A(net151741), .Y(net147506) );
  INVX1 U8846 ( .A(n20943), .Y(n20942) );
  INVX1 U8847 ( .A(net142728), .Y(n20943) );
  AOI22X1 U8848 ( .A(n4199), .B(net151751), .C(n3285), .D(n20942), .Y(net90010) );
  BUFX2 U8849 ( .A(n20944), .Y(net142728) );
  INVX1 U8850 ( .A(n20943), .Y(net151649) );
  INVX1 U8851 ( .A(net107076), .Y(net107094) );
  AOI21X1 U8852 ( .A(n20946), .B(n20950), .C(reset), .Y(n20944) );
  BUFX2 U8853 ( .A(n20951), .Y(n20946) );
  NAND3X1 U8854 ( .A(net95147), .B(net103869), .C(net147735), .Y(n20951) );
  AND2X2 U8855 ( .A(net109585), .B(net125066), .Y(net95147) );
  BUFX2 U8856 ( .A(net90052), .Y(net103869) );
  AND2X2 U8857 ( .A(net111600), .B(n14346), .Y(n20950) );
  INVX1 U8858 ( .A(net90053), .Y(net111600) );
  INVX1 U8859 ( .A(net114546), .Y(n14346) );
  INVX1 U8860 ( .A(n34242), .Y(n20952) );
  MUX2X1 U8861 ( .B(grid[382]), .A(grid[376]), .S(net105778), .Y(n28162) );
  BUFX2 U8862 ( .A(net110927), .Y(net151977) );
  AND2X2 U8863 ( .A(n21135), .B(n25467), .Y(n21322) );
  INVX1 U8864 ( .A(n20973), .Y(n20953) );
  INVX2 U8865 ( .A(n34443), .Y(n25621) );
  INVX1 U8866 ( .A(n25649), .Y(n25636) );
  INVX1 U8867 ( .A(n25727), .Y(n20954) );
  INVX1 U8868 ( .A(n20954), .Y(n20955) );
  AND2X2 U8869 ( .A(n33052), .B(n33051), .Y(n20956) );
  INVX2 U8870 ( .A(net116754), .Y(net151617) );
  MUX2X1 U8871 ( .B(grid[304]), .A(grid[310]), .S(net150251), .Y(n28171) );
  MUX2X1 U8872 ( .B(grid[16]), .A(grid[22]), .S(net112202), .Y(n28216) );
  INVX1 U8873 ( .A(net111984), .Y(net151886) );
  INVX1 U8874 ( .A(net151886), .Y(net151887) );
  MUX2X1 U8875 ( .B(n28020), .A(n28035), .S(net89785), .Y(n28038) );
  INVX1 U8876 ( .A(n29369), .Y(n20966) );
  INVX1 U8877 ( .A(n29369), .Y(n20957) );
  INVX1 U8878 ( .A(n29369), .Y(n20958) );
  INVX1 U8879 ( .A(net151709), .Y(net151875) );
  BUFX2 U8880 ( .A(n33905), .Y(n20959) );
  INVX2 U8881 ( .A(n11049), .Y(n21240) );
  XOR2X1 U8882 ( .A(n34312), .B(n20960), .Y(n34314) );
  XNOR2X1 U8883 ( .A(n23203), .B(n34317), .Y(n20960) );
  INVX1 U8884 ( .A(net107074), .Y(net151840) );
  INVX1 U8885 ( .A(n20974), .Y(n20961) );
  BUFX2 U8886 ( .A(alt14_net96296), .Y(net151833) );
  BUFX2 U8887 ( .A(alt14_net96296), .Y(net151834) );
  INVX1 U8888 ( .A(n25649), .Y(n25650) );
  INVX1 U8889 ( .A(n29369), .Y(n23209) );
  INVX1 U8890 ( .A(net151812), .Y(net107061) );
  INVX1 U8891 ( .A(net112181), .Y(net151814) );
  INVX1 U8892 ( .A(net142728), .Y(net151812) );
  AND2X2 U8893 ( .A(n22048), .B(n23927), .Y(n21840) );
  INVX2 U8894 ( .A(n11047), .Y(n21241) );
  MUX2X1 U8895 ( .B(grid[320]), .A(grid[314]), .S(net116777), .Y(n28047) );
  INVX1 U8896 ( .A(net149909), .Y(net151801) );
  BUFX2 U8897 ( .A(n3244), .Y(n20962) );
  BUFX2 U8898 ( .A(n34270), .Y(n20963) );
  NOR3X1 U8899 ( .A(n20965), .B(n21148), .C(n34327), .Y(n20964) );
  INVX8 U8900 ( .A(n34328), .Y(n20965) );
  OR2X2 U8901 ( .A(n29369), .B(n34134), .Y(n21744) );
  OR2X2 U8902 ( .A(n29369), .B(n34135), .Y(n21745) );
  OR2X2 U8903 ( .A(n29369), .B(n34136), .Y(n21746) );
  OR2X2 U8904 ( .A(n29369), .B(n34137), .Y(n21747) );
  OR2X2 U8905 ( .A(n29369), .B(n34138), .Y(n21748) );
  OR2X2 U8906 ( .A(n29369), .B(n34139), .Y(n21749) );
  OR2X2 U8907 ( .A(n29369), .B(n34140), .Y(n21750) );
  OR2X2 U8908 ( .A(n29369), .B(n34141), .Y(n21751) );
  OR2X2 U8909 ( .A(n29369), .B(n34142), .Y(n21752) );
  OR2X2 U8910 ( .A(n29369), .B(n34143), .Y(n21753) );
  OR2X2 U8911 ( .A(n29369), .B(n34144), .Y(n21754) );
  OR2X2 U8912 ( .A(n29369), .B(n34145), .Y(n21755) );
  INVX4 U8913 ( .A(n21161), .Y(n29369) );
  AND2X2 U8914 ( .A(n34350), .B(n25588), .Y(n34373) );
  OR2X2 U8915 ( .A(n34281), .B(n25662), .Y(n11047) );
  INVX1 U8916 ( .A(net151741), .Y(net151751) );
  INVX1 U8917 ( .A(net147481), .Y(net151741) );
  INVX1 U8918 ( .A(net151741), .Y(net151738) );
  INVX1 U8919 ( .A(n25728), .Y(n20967) );
  INVX1 U8920 ( .A(n25728), .Y(n34380) );
  INVX2 U8921 ( .A(n34244), .Y(n34242) );
  AND2X1 U8922 ( .A(net95147), .B(net96340), .Y(n25482) );
  INVX4 U8923 ( .A(n25482), .Y(n29383) );
  INVX1 U8924 ( .A(net151709), .Y(net151710) );
  INVX1 U8925 ( .A(net151629), .Y(net151696) );
  INVX1 U8926 ( .A(net151629), .Y(net151697) );
  INVX1 U8927 ( .A(net151629), .Y(net116760) );
  INVX4 U8928 ( .A(n29606), .Y(n20968) );
  INVX2 U8929 ( .A(oc[18]), .Y(n29606) );
  BUFX2 U8930 ( .A(n34441), .Y(n20969) );
  INVX1 U8931 ( .A(n25851), .Y(n20970) );
  INVX4 U8932 ( .A(n29193), .Y(n34441) );
  INVX1 U8933 ( .A(net111237), .Y(net151662) );
  INVX1 U8934 ( .A(net151633), .Y(net151652) );
  MUX2X1 U8935 ( .B(n28081), .A(n28080), .S(net105822), .Y(n28079) );
  INVX2 U8936 ( .A(net105810), .Y(net105822) );
  MUX2X1 U8937 ( .B(n28045), .A(n28044), .S(net105822), .Y(n28043) );
  INVX1 U8938 ( .A(net109766), .Y(net151632) );
  INVX1 U8939 ( .A(net151632), .Y(net151633) );
  INVX1 U8940 ( .A(net151662), .Y(net151629) );
  MUX2X1 U8941 ( .B(n28084), .A(n28083), .S(net151626), .Y(n28082) );
  INVX8 U8942 ( .A(net113954), .Y(net151626) );
  XNOR2X1 U8943 ( .A(n34433), .B(n34432), .Y(n34435) );
  INVX1 U8944 ( .A(n22676), .Y(n20971) );
  INVX1 U8945 ( .A(n29527), .Y(n20972) );
  XNOR2X1 U8946 ( .A(n34234), .B(n34441), .Y(n20973) );
  INVX1 U8947 ( .A(n20973), .Y(n34235) );
  AND2X2 U8948 ( .A(n22085), .B(n34267), .Y(n34269) );
  OR2X2 U8949 ( .A(oc[20]), .B(oc[22]), .Y(n29607) );
  INVX1 U8950 ( .A(n3774), .Y(n34279) );
  INVX1 U8951 ( .A(n33078), .Y(n33077) );
  BUFX2 U8952 ( .A(n26168), .Y(n26175) );
  BUFX2 U8953 ( .A(n26169), .Y(n26176) );
  BUFX2 U8954 ( .A(n26171), .Y(n26178) );
  BUFX2 U8955 ( .A(n26170), .Y(n26177) );
  INVX2 U8956 ( .A(oc[5]), .Y(n29946) );
  INVX2 U8957 ( .A(n26338), .Y(n30186) );
  INVX1 U8958 ( .A(n33105), .Y(n33145) );
  INVX1 U8959 ( .A(n34421), .Y(n21108) );
  INVX1 U8960 ( .A(n25069), .Y(n21111) );
  AND2X1 U8961 ( .A(n27076), .B(n27000), .Y(n16026) );
  AND2X1 U8962 ( .A(n26867), .B(n26933), .Y(n16103) );
  AND2X1 U8963 ( .A(n26929), .B(n27086), .Y(n16184) );
  AND2X1 U8964 ( .A(n26995), .B(n27177), .Y(n15952) );
  AND2X1 U8965 ( .A(n26918), .B(n26857), .Y(n16010) );
  AND2X1 U8966 ( .A(n25341), .B(n24940), .Y(n16083) );
  AND2X1 U8967 ( .A(n25151), .B(n25156), .Y(n16087) );
  OR2X1 U8968 ( .A(n27077), .B(n16114), .Y(n16121) );
  AND2X1 U8969 ( .A(n23594), .B(n23741), .Y(n16088) );
  OR2X1 U8970 ( .A(n27086), .B(n16211), .Y(n16219) );
  AND2X1 U8971 ( .A(n26918), .B(n26804), .Y(n16163) );
  AND2X1 U8972 ( .A(n26805), .B(n26938), .Y(n16158) );
  OR2X1 U8973 ( .A(n27177), .B(n15979), .Y(n15987) );
  AND2X1 U8974 ( .A(n26999), .B(n24942), .Y(n15932) );
  AND2X1 U8975 ( .A(n26917), .B(n25157), .Y(n15936) );
  INVX1 U8976 ( .A(n21126), .Y(n33061) );
  INVX1 U8977 ( .A(n32476), .Y(n25745) );
  AND2X1 U8978 ( .A(n23595), .B(n23742), .Y(n16011) );
  OR2X1 U8979 ( .A(n27193), .B(n16195), .Y(n16044) );
  AND2X1 U8980 ( .A(n23641), .B(n25198), .Y(n16092) );
  OR2X1 U8981 ( .A(n34579), .B(n27183), .Y(n16098) );
  AND2X1 U8982 ( .A(n23593), .B(n23740), .Y(n16169) );
  OR2X1 U8983 ( .A(n27193), .B(n16195), .Y(n16202) );
  AND2X1 U8984 ( .A(n26858), .B(n26918), .Y(n16166) );
  AND2X1 U8985 ( .A(n29649), .B(n27113), .Y(n27274) );
  OR2X1 U8986 ( .A(n26930), .B(n15963), .Y(n15970) );
  AND2X1 U8987 ( .A(n23596), .B(n23743), .Y(n15937) );
  INVX1 U8988 ( .A(n26491), .Y(n21075) );
  INVX1 U8989 ( .A(n21146), .Y(n21235) );
  INVX1 U8990 ( .A(n25604), .Y(n34353) );
  AND2X1 U8991 ( .A(n23642), .B(n25200), .Y(n15941) );
  INVX1 U8992 ( .A(n28608), .Y(n21077) );
  INVX1 U8993 ( .A(n28607), .Y(n21079) );
  AND2X1 U8994 ( .A(n26897), .B(n29614), .Y(n29616) );
  INVX1 U8995 ( .A(n25585), .Y(n34293) );
  INVX2 U8996 ( .A(n34402), .Y(n34390) );
  INVX1 U8997 ( .A(n29486), .Y(n21032) );
  INVX1 U8998 ( .A(n27172), .Y(n21170) );
  AND2X1 U8999 ( .A(n32607), .B(n32608), .Y(n32609) );
  INVX1 U9000 ( .A(n34410), .Y(n21148) );
  OR2X1 U9001 ( .A(n24016), .B(n24018), .Y(n29691) );
  OR2X1 U9002 ( .A(n30076), .B(n29320), .Y(n30077) );
  AND2X1 U9003 ( .A(n25164), .B(n25468), .Y(n25469) );
  INVX1 U9004 ( .A(n25411), .Y(n29252) );
  INVX2 U9005 ( .A(n29266), .Y(n21006) );
  INVX2 U9006 ( .A(n25698), .Y(n25756) );
  AND2X1 U9007 ( .A(n29730), .B(n27018), .Y(n27248) );
  INVX1 U9008 ( .A(loc_s2[4]), .Y(n21208) );
  INVX1 U9009 ( .A(n33147), .Y(n33142) );
  INVX1 U9010 ( .A(n25435), .Y(n34307) );
  INVX1 U9011 ( .A(n23277), .Y(n34432) );
  OR2X1 U9012 ( .A(n27192), .B(n29469), .Y(n14478) );
  AND2X1 U9013 ( .A(n29525), .B(n29524), .Y(n32185) );
  AND2X1 U9014 ( .A(n22950), .B(n27018), .Y(n27249) );
  INVX1 U9015 ( .A(direction_line[0]), .Y(n21238) );
  AND2X1 U9016 ( .A(n23590), .B(n25841), .Y(n29696) );
  OR2X1 U9017 ( .A(n20975), .B(n27192), .Y(n14871) );
  AND2X1 U9018 ( .A(n23643), .B(n30479), .Y(n30484) );
  OR2X1 U9019 ( .A(n31649), .B(n31650), .Y(n31651) );
  AND2X1 U9020 ( .A(n34174), .B(net103869), .Y(n32198) );
  INVX1 U9021 ( .A(n27159), .Y(n21128) );
  INVX1 U9022 ( .A(n33450), .Y(n21065) );
  INVX1 U9023 ( .A(n12020), .Y(n21064) );
  INVX1 U9024 ( .A(n33467), .Y(n21062) );
  INVX1 U9025 ( .A(n12015), .Y(n21061) );
  INVX1 U9026 ( .A(n33473), .Y(n21053) );
  INVX1 U9027 ( .A(n12014), .Y(n21052) );
  AND2X1 U9028 ( .A(n24943), .B(n30021), .Y(n29881) );
  INVX1 U9029 ( .A(n33614), .Y(n21050) );
  INVX1 U9030 ( .A(n11979), .Y(n21049) );
  AND2X1 U9031 ( .A(n30038), .B(n26982), .Y(n29767) );
  AND2X1 U9032 ( .A(n23479), .B(n25107), .Y(n29753) );
  INVX1 U9033 ( .A(n25408), .Y(n29565) );
  INVX1 U9034 ( .A(n26485), .Y(n26515) );
  AND2X1 U9035 ( .A(n27273), .B(n27114), .Y(n30027) );
  INVX1 U9036 ( .A(n25344), .Y(n25458) );
  AND2X1 U9037 ( .A(n23591), .B(n21432), .Y(n15897) );
  AND2X1 U9038 ( .A(n23480), .B(n23649), .Y(n15156) );
  AND2X1 U9039 ( .A(n23481), .B(n23650), .Y(n15143) );
  AND2X1 U9040 ( .A(n23482), .B(n23651), .Y(n15131) );
  AND2X1 U9041 ( .A(n23483), .B(n23652), .Y(n15119) );
  AND2X1 U9042 ( .A(n23484), .B(n23653), .Y(n15107) );
  AND2X1 U9043 ( .A(n23485), .B(n23654), .Y(n15095) );
  AND2X1 U9044 ( .A(n23486), .B(n23655), .Y(n15083) );
  AND2X1 U9045 ( .A(n23487), .B(n23656), .Y(n15071) );
  AND2X1 U9046 ( .A(n23488), .B(n23657), .Y(n15058) );
  AND2X1 U9047 ( .A(n23489), .B(n23658), .Y(n15046) );
  AND2X1 U9048 ( .A(n23490), .B(n23659), .Y(n15034) );
  AND2X1 U9049 ( .A(n23491), .B(n23660), .Y(n15022) );
  AND2X1 U9050 ( .A(n23492), .B(n23661), .Y(n15010) );
  AND2X1 U9051 ( .A(n23493), .B(n23662), .Y(n14998) );
  AND2X1 U9052 ( .A(n23494), .B(n23663), .Y(n14986) );
  AND2X1 U9053 ( .A(n23495), .B(n23664), .Y(n14974) );
  AND2X1 U9054 ( .A(n23496), .B(n23665), .Y(n14960) );
  AND2X1 U9055 ( .A(n23497), .B(n23666), .Y(n14948) );
  AND2X1 U9056 ( .A(n23498), .B(n23667), .Y(n14936) );
  AND2X1 U9057 ( .A(n23499), .B(n23668), .Y(n14924) );
  AND2X1 U9058 ( .A(n23500), .B(n23669), .Y(n14912) );
  AND2X1 U9059 ( .A(n23501), .B(n23670), .Y(n14900) );
  AND2X1 U9060 ( .A(n23502), .B(n23671), .Y(n14888) );
  AND2X1 U9061 ( .A(n23503), .B(n23672), .Y(n14876) );
  AND2X1 U9062 ( .A(n23504), .B(n23673), .Y(n14862) );
  AND2X1 U9063 ( .A(n23505), .B(n23674), .Y(n14850) );
  AND2X1 U9064 ( .A(n23506), .B(n23675), .Y(n14838) );
  AND2X1 U9065 ( .A(n23507), .B(n23676), .Y(n14826) );
  AND2X1 U9066 ( .A(n23508), .B(n23677), .Y(n14814) );
  AND2X1 U9067 ( .A(n23509), .B(n23678), .Y(n14802) );
  AND2X1 U9068 ( .A(n23510), .B(n23679), .Y(n14790) );
  AND2X1 U9069 ( .A(n23511), .B(n23680), .Y(n14778) );
  AND2X1 U9070 ( .A(n23512), .B(n23681), .Y(n14764) );
  AND2X1 U9071 ( .A(n23513), .B(n23682), .Y(n14752) );
  AND2X1 U9072 ( .A(n23514), .B(n23683), .Y(n14740) );
  AND2X1 U9073 ( .A(n23515), .B(n23684), .Y(n14728) );
  AND2X1 U9074 ( .A(n23516), .B(n23685), .Y(n14716) );
  AND2X1 U9075 ( .A(n23517), .B(n23686), .Y(n14704) );
  AND2X1 U9076 ( .A(n23518), .B(n23687), .Y(n14692) );
  AND2X1 U9077 ( .A(n23519), .B(n23688), .Y(n14680) );
  AND2X1 U9078 ( .A(n23520), .B(n23689), .Y(n14665) );
  AND2X1 U9079 ( .A(n23521), .B(n23690), .Y(n14653) );
  AND2X1 U9080 ( .A(n23522), .B(n23691), .Y(n14641) );
  AND2X1 U9081 ( .A(n23523), .B(n23692), .Y(n14629) );
  AND2X1 U9082 ( .A(n23524), .B(n23693), .Y(n14617) );
  AND2X1 U9083 ( .A(n23525), .B(n23694), .Y(n14605) );
  AND2X1 U9084 ( .A(n23526), .B(n23695), .Y(n14593) );
  AND2X1 U9085 ( .A(n23527), .B(n23696), .Y(n14581) );
  AND2X1 U9086 ( .A(n23528), .B(n23697), .Y(n14567) );
  AND2X1 U9087 ( .A(n23529), .B(n23698), .Y(n14555) );
  AND2X1 U9088 ( .A(n23530), .B(n23699), .Y(n14543) );
  AND2X1 U9089 ( .A(n23531), .B(n23700), .Y(n14531) );
  AND2X1 U9090 ( .A(n23532), .B(n23701), .Y(n14519) );
  AND2X1 U9091 ( .A(n23533), .B(n23702), .Y(n14507) );
  AND2X1 U9092 ( .A(n23534), .B(n23703), .Y(n14495) );
  AND2X1 U9093 ( .A(n23535), .B(n23704), .Y(n14483) );
  AND2X1 U9094 ( .A(n23536), .B(n23705), .Y(n14468) );
  AND2X1 U9095 ( .A(n23537), .B(n23706), .Y(n14455) );
  AND2X1 U9096 ( .A(n23538), .B(n23707), .Y(n14442) );
  AND2X1 U9097 ( .A(n23539), .B(n23708), .Y(n14429) );
  AND2X1 U9098 ( .A(n23540), .B(n23709), .Y(n14416) );
  AND2X1 U9099 ( .A(n23541), .B(n23710), .Y(n14403) );
  AND2X1 U9100 ( .A(n23542), .B(n23711), .Y(n14390) );
  OR2X1 U9101 ( .A(n24017), .B(n30483), .Y(n14372) );
  AND2X1 U9102 ( .A(n23589), .B(n23647), .Y(n16269) );
  AND2X1 U9103 ( .A(n23592), .B(n23648), .Y(n15245) );
  AND2X1 U9104 ( .A(n21543), .B(n23744), .Y(n34487) );
  INVX1 U9105 ( .A(n21839), .Y(n21293) );
  INVX1 U9106 ( .A(n21829), .Y(n21302) );
  INVX1 U9107 ( .A(n21826), .Y(n21305) );
  INVX1 U9108 ( .A(n21823), .Y(n23626) );
  AND2X1 U9109 ( .A(n21533), .B(n23939), .Y(n21823) );
  INVX1 U9110 ( .A(n21821), .Y(n21308) );
  AND2X1 U9111 ( .A(n23478), .B(n29733), .Y(n15887) );
  INVX1 U9112 ( .A(n21854), .Y(n21354) );
  INVX1 U9113 ( .A(n25829), .Y(n21846) );
  AND2X1 U9114 ( .A(n21540), .B(n23746), .Y(n25829) );
  INVX1 U9115 ( .A(n21107), .Y(n34440) );
  INVX1 U9116 ( .A(n21832), .Y(n21299) );
  AND2X2 U9117 ( .A(n22052), .B(n23931), .Y(n21832) );
  INVX1 U9118 ( .A(n20956), .Y(n20974) );
  INVX2 U9119 ( .A(n20961), .Y(n25649) );
  BUFX2 U9120 ( .A(n25620), .Y(n27917) );
  INVX8 U9121 ( .A(n25441), .Y(n33308) );
  INVX2 U9122 ( .A(n33002), .Y(n25441) );
  INVX2 U9123 ( .A(n2245), .Y(n28987) );
  INVX1 U9124 ( .A(n27223), .Y(n29442) );
  INVX8 U9125 ( .A(n29282), .Y(n29277) );
  INVX8 U9126 ( .A(n29419), .Y(n29414) );
  AND2X1 U9127 ( .A(T[3]), .B(n24941), .Y(n34574) );
  INVX4 U9128 ( .A(n20809), .Y(n21066) );
  AND2X1 U9129 ( .A(n24937), .B(n34360), .Y(n16104) );
  AND2X1 U9130 ( .A(n25109), .B(n34385), .Y(n16122) );
  INVX8 U9131 ( .A(n23107), .Y(n21106) );
  AND2X1 U9132 ( .A(n21545), .B(n21423), .Y(n27140) );
  AND2X1 U9133 ( .A(n21526), .B(n23646), .Y(net89759) );
  INVX1 U9134 ( .A(n29404), .Y(n29403) );
  INVX1 U9135 ( .A(n29421), .Y(n29420) );
  INVX1 U9136 ( .A(n29413), .Y(n29412) );
  AND2X1 U9137 ( .A(n26753), .B(n26871), .Y(n29642) );
  AND2X1 U9138 ( .A(n34210), .B(n29476), .Y(n29481) );
  INVX1 U9139 ( .A(n23274), .Y(n26978) );
  AND2X1 U9140 ( .A(n30673), .B(net96340), .Y(n30687) );
  AND2X1 U9141 ( .A(n30855), .B(net96340), .Y(n30866) );
  AND2X1 U9142 ( .A(n31014), .B(net96340), .Y(n31025) );
  AND2X1 U9143 ( .A(n31092), .B(net96340), .Y(n31103) );
  AND2X1 U9144 ( .A(n31560), .B(net96340), .Y(n31571) );
  INVX8 U9145 ( .A(n29464), .Y(n28599) );
  AND2X1 U9146 ( .A(n31502), .B(net96340), .Y(n31512) );
  INVX8 U9147 ( .A(n26764), .Y(n26077) );
  INVX1 U9148 ( .A(n24936), .Y(n21408) );
  INVX8 U9149 ( .A(n8053), .Y(n29461) );
  INVX1 U9150 ( .A(n26260), .Y(n26268) );
  INVX2 U9151 ( .A(n33019), .Y(n26078) );
  BUFX2 U9152 ( .A(n27147), .Y(n29212) );
  INVX2 U9153 ( .A(n29465), .Y(n29185) );
  AND2X1 U9154 ( .A(n29221), .B(n26793), .Y(n30683) );
  AND2X1 U9155 ( .A(n29221), .B(n26861), .Y(n30706) );
  AND2X1 U9156 ( .A(n29221), .B(n26746), .Y(n30726) );
  AND2X1 U9157 ( .A(n29221), .B(n26706), .Y(n30766) );
  AND2X1 U9158 ( .A(n29221), .B(n26675), .Y(n30806) );
  AND2X1 U9159 ( .A(n29221), .B(n24945), .Y(n30846) );
  AND2X1 U9160 ( .A(n29221), .B(n24946), .Y(n30886) );
  AND2X1 U9161 ( .A(n29221), .B(n26921), .Y(n30906) );
  AND2X1 U9162 ( .A(n29221), .B(n26847), .Y(n30927) );
  AND2X1 U9163 ( .A(n29221), .B(n26792), .Y(n30967) );
  AND2X1 U9164 ( .A(n29221), .B(n26791), .Y(n30987) );
  AND2X1 U9165 ( .A(n29221), .B(n26745), .Y(n31024) );
  AND2X1 U9166 ( .A(n29221), .B(n24947), .Y(n31062) );
  AND2X1 U9167 ( .A(n29221), .B(n24948), .Y(n31102) );
  AND2X1 U9168 ( .A(n29221), .B(n24949), .Y(n31142) );
  AND2X1 U9169 ( .A(n29221), .B(n24950), .Y(n31179) );
  AND2X1 U9170 ( .A(n29221), .B(n24951), .Y(n31219) );
  AND2X1 U9171 ( .A(n29221), .B(n24952), .Y(n31259) );
  AND2X1 U9172 ( .A(n29221), .B(n26860), .Y(n31296) );
  AND2X1 U9173 ( .A(n29221), .B(n26744), .Y(n31315) );
  AND2X1 U9174 ( .A(n29221), .B(n26790), .Y(n31353) );
  AND2X1 U9175 ( .A(n29221), .B(n26674), .Y(n31393) );
  AND2X1 U9176 ( .A(n29221), .B(n24953), .Y(n31434) );
  AND2X1 U9177 ( .A(n29221), .B(n24954), .Y(n31473) );
  AND2X1 U9178 ( .A(n29221), .B(n24955), .Y(n31511) );
  AND2X1 U9179 ( .A(n29221), .B(n27066), .Y(n31530) );
  AND2X1 U9180 ( .A(n29221), .B(n26789), .Y(n31550) );
  AND2X1 U9181 ( .A(n29221), .B(n26846), .Y(n31591) );
  AND2X1 U9182 ( .A(n29221), .B(n26743), .Y(n31610) );
  AND2X1 U9183 ( .A(n29221), .B(n26705), .Y(n31646) );
  AND2X1 U9184 ( .A(n29221), .B(n24956), .Y(n31685) );
  AND2X1 U9185 ( .A(n29221), .B(n24957), .Y(n31724) );
  AND2X1 U9186 ( .A(n29221), .B(n24958), .Y(n31762) );
  AND2X1 U9187 ( .A(n29221), .B(n24959), .Y(n31802) );
  AND2X1 U9188 ( .A(n29221), .B(n24960), .Y(n31841) );
  AND2X1 U9189 ( .A(n29221), .B(n24961), .Y(n31882) );
  AND2X1 U9190 ( .A(n24938), .B(n34360), .Y(n16027) );
  AND2X1 U9191 ( .A(n27273), .B(n26981), .Y(n30496) );
  INVX1 U9192 ( .A(n33993), .Y(n21204) );
  AND2X1 U9193 ( .A(n21432), .B(n22990), .Y(n27273) );
  INVX1 U9194 ( .A(n34616), .Y(n20975) );
  INVX1 U9195 ( .A(address[1]), .Y(n29471) );
  INVX1 U9196 ( .A(address[2]), .Y(n29470) );
  INVX1 U9197 ( .A(net114916), .Y(net151429) );
  INVX1 U9198 ( .A(net113955), .Y(net114916) );
  INVX1 U9199 ( .A(n28220), .Y(n21130) );
  BUFX2 U9200 ( .A(n32166), .Y(n20976) );
  AND2X1 U9201 ( .A(n29592), .B(n29591), .Y(n29596) );
  INVX1 U9202 ( .A(n29582), .Y(n29592) );
  INVX1 U9203 ( .A(n21203), .Y(n20977) );
  INVX1 U9204 ( .A(n21203), .Y(n21184) );
  INVX1 U9205 ( .A(n21325), .Y(n26949) );
  OR2X2 U9206 ( .A(n33934), .B(reset), .Y(n21325) );
  BUFX2 U9207 ( .A(address[0]), .Y(n20978) );
  INVX2 U9208 ( .A(n23276), .Y(n25346) );
  INVX1 U9209 ( .A(n20991), .Y(n20979) );
  INVX1 U9210 ( .A(n31921), .Y(n20980) );
  INVX1 U9211 ( .A(n31921), .Y(n20981) );
  INVX1 U9212 ( .A(n20991), .Y(n20982) );
  INVX1 U9213 ( .A(n20993), .Y(n20983) );
  INVX1 U9214 ( .A(n20982), .Y(n20984) );
  INVX1 U9215 ( .A(n20982), .Y(n20985) );
  INVX1 U9216 ( .A(n20988), .Y(n20986) );
  INVX1 U9217 ( .A(n31921), .Y(n20987) );
  INVX1 U9218 ( .A(n20991), .Y(n20988) );
  INVX1 U9219 ( .A(n20992), .Y(n20989) );
  INVX2 U9220 ( .A(n29313), .Y(n25740) );
  INVX1 U9221 ( .A(n20979), .Y(n20990) );
  AND2X2 U9222 ( .A(n20995), .B(n27152), .Y(n20991) );
  INVX1 U9223 ( .A(n27224), .Y(n20992) );
  INVX1 U9224 ( .A(n20991), .Y(n20993) );
  INVX1 U9225 ( .A(n27173), .Y(n20994) );
  INVX1 U9226 ( .A(n27173), .Y(n34196) );
  OR2X2 U9227 ( .A(n22102), .B(n27157), .Y(n20995) );
  AND2X2 U9228 ( .A(n20995), .B(n27152), .Y(n20996) );
  AND2X2 U9229 ( .A(net96340), .B(n31675), .Y(n31686) );
  INVX1 U9230 ( .A(n25694), .Y(n20534) );
  INVX8 U9231 ( .A(n31891), .Y(n26324) );
  AND2X2 U9232 ( .A(net96340), .B(n31792), .Y(n31803) );
  AND2X2 U9233 ( .A(n30696), .B(net96340), .Y(n30707) );
  INVX1 U9234 ( .A(n29209), .Y(n20997) );
  INVX1 U9235 ( .A(n34209), .Y(n20998) );
  INVX1 U9236 ( .A(n20998), .Y(n20999) );
  INVX1 U9237 ( .A(n25411), .Y(n21000) );
  INVX1 U9238 ( .A(n29236), .Y(n21001) );
  INVX1 U9239 ( .A(n29236), .Y(n21002) );
  INVX1 U9240 ( .A(n29236), .Y(n21003) );
  INVX1 U9241 ( .A(n29236), .Y(n29232) );
  INVX1 U9242 ( .A(n26463), .Y(n21004) );
  INVX1 U9243 ( .A(net114723), .Y(net151212) );
  INVX1 U9244 ( .A(n21404), .Y(n21271) );
  XOR2X1 U9245 ( .A(alt5_net95668), .B(n2252), .Y(n21156) );
  MUX2X1 U9246 ( .B(n29595), .A(n34503), .S(n21156), .Y(n29562) );
  OAI21X1 U9247 ( .A(n21006), .B(n23422), .C(n26294), .Y(n21005) );
  INVX1 U9248 ( .A(n21005), .Y(n31869) );
  AND2X2 U9249 ( .A(n27257), .B(n23441), .Y(n27307) );
  AND2X2 U9250 ( .A(n29683), .B(n30127), .Y(n27257) );
  INVX1 U9251 ( .A(n30127), .Y(n21007) );
  AND2X2 U9252 ( .A(net96340), .B(n31323), .Y(n31334) );
  OAI21X1 U9253 ( .A(n29271), .B(n23373), .C(n26286), .Y(n21008) );
  INVX1 U9254 ( .A(n21008), .Y(n31422) );
  OAI21X1 U9255 ( .A(n29271), .B(n23365), .C(n26286), .Y(n21009) );
  INVX1 U9256 ( .A(n21009), .Y(n31341) );
  OR2X2 U9257 ( .A(n23254), .B(n31504), .Y(n21010) );
  INVX1 U9258 ( .A(n34612), .Y(n21011) );
  INVX1 U9259 ( .A(n29488), .Y(n21012) );
  AND2X2 U9260 ( .A(n21069), .B(n21557), .Y(n21013) );
  OR2X2 U9261 ( .A(n23261), .B(n31563), .Y(n21014) );
  OR2X2 U9262 ( .A(n23268), .B(n31717), .Y(n21015) );
  OR2X2 U9263 ( .A(n23213), .B(n30676), .Y(n21016) );
  OR2X2 U9264 ( .A(n23239), .B(n30858), .Y(n21017) );
  OR2X2 U9265 ( .A(n23622), .B(n31017), .Y(n21018) );
  OR2X2 U9266 ( .A(n23625), .B(n31584), .Y(n21019) );
  OAI21X1 U9267 ( .A(n29271), .B(n23336), .C(n26295), .Y(n21020) );
  INVX1 U9268 ( .A(n21020), .Y(n31050) );
  OR2X2 U9269 ( .A(n23216), .B(n30699), .Y(n21021) );
  OAI21X1 U9270 ( .A(n29271), .B(n32000), .C(n26281), .Y(n21022) );
  INVX1 U9271 ( .A(n21022), .Y(n30996) );
  INVX1 U9272 ( .A(n21011), .Y(n21023) );
  INVX1 U9273 ( .A(n22674), .Y(n21024) );
  INVX1 U9274 ( .A(n22674), .Y(n29490) );
  OR2X2 U9275 ( .A(n23219), .B(n30719), .Y(n21025) );
  OR2X2 U9276 ( .A(n23251), .B(n31252), .Y(n21026) );
  OAI21X1 U9277 ( .A(n29270), .B(n23360), .C(n26288), .Y(n21027) );
  INVX1 U9278 ( .A(n21027), .Y(n31304) );
  OR2X2 U9279 ( .A(n29487), .B(n21032), .Y(n21028) );
  INVX1 U9280 ( .A(n25570), .Y(n21029) );
  BUFX2 U9281 ( .A(locTrig[0]), .Y(n21030) );
  INVX4 U9282 ( .A(n27906), .Y(n33062) );
  OR2X2 U9283 ( .A(n29487), .B(n21032), .Y(n21031) );
  INVX1 U9284 ( .A(n25674), .Y(n21033) );
  OR2X2 U9285 ( .A(n23242), .B(n30920), .Y(n21034) );
  OR2X2 U9286 ( .A(n23248), .B(n31212), .Y(n21035) );
  OR2X2 U9287 ( .A(n23229), .B(n30778), .Y(n21036) );
  BUFX4 U9288 ( .A(n29204), .Y(n29197) );
  OAI21X1 U9289 ( .A(n29271), .B(n23413), .C(n26294), .Y(n21037) );
  INVX1 U9290 ( .A(n21037), .Y(n31790) );
  INVX4 U9291 ( .A(n29271), .Y(n29266) );
  INVX1 U9292 ( .A(n30867), .Y(n21038) );
  OAI21X1 U9293 ( .A(n29271), .B(n31978), .C(n26294), .Y(n21039) );
  INVX1 U9294 ( .A(n21039), .Y(n30894) );
  INVX1 U9295 ( .A(n30728), .Y(n21040) );
  OR2X2 U9296 ( .A(n23235), .B(n21041), .Y(n23234) );
  OR2X2 U9297 ( .A(n23236), .B(n30818), .Y(n21041) );
  AND2X2 U9298 ( .A(n29289), .B(n31909), .Y(n21042) );
  INVX2 U9299 ( .A(n29289), .Y(n29287) );
  INVX1 U9300 ( .A(n26514), .Y(n21043) );
  INVX8 U9301 ( .A(n21096), .Y(n26514) );
  AND2X2 U9302 ( .A(n22983), .B(n22995), .Y(n21044) );
  OAI21X1 U9303 ( .A(n29270), .B(n31943), .C(n26288), .Y(n21045) );
  INVX1 U9304 ( .A(n21045), .Y(n30754) );
  INVX1 U9305 ( .A(n29270), .Y(n29269) );
  INVX1 U9306 ( .A(n30929), .Y(n21046) );
  INVX1 U9307 ( .A(n30747), .Y(n21047) );
  OAI21X1 U9308 ( .A(n21049), .B(net96596), .C(n21050), .Y(n21048) );
  INVX1 U9309 ( .A(n21048), .Y(n33616) );
  OAI21X1 U9310 ( .A(n21052), .B(net96596), .C(n21053), .Y(n21051) );
  INVX1 U9311 ( .A(n21051), .Y(n33475) );
  OAI21X1 U9312 ( .A(n29271), .B(n23390), .C(n26294), .Y(n21054) );
  INVX1 U9313 ( .A(n21054), .Y(n31579) );
  INVX2 U9314 ( .A(n29271), .Y(n29267) );
  INVX2 U9315 ( .A(n29477), .Y(n27084) );
  INVX1 U9316 ( .A(n27019), .Y(n21055) );
  INVX1 U9317 ( .A(n26278), .Y(n26293) );
  INVX1 U9318 ( .A(n26295), .Y(n21056) );
  INVX1 U9319 ( .A(n30073), .Y(n21057) );
  INVX2 U9320 ( .A(n26514), .Y(n26500) );
  INVX1 U9321 ( .A(n30638), .Y(n21058) );
  INVX1 U9322 ( .A(n21192), .Y(n21059) );
  MUX2X1 U9323 ( .B(n28237), .A(n28240), .S(n28602), .Y(n28251) );
  OAI21X1 U9324 ( .A(n21061), .B(net96596), .C(n21062), .Y(n21060) );
  INVX1 U9325 ( .A(n21060), .Y(n33469) );
  OAI21X1 U9326 ( .A(n21064), .B(net96596), .C(n21065), .Y(n21063) );
  INVX1 U9327 ( .A(n21063), .Y(n33452) );
  MUX2X1 U9328 ( .B(n28577), .A(n28580), .S(n21066), .Y(n28591) );
  INVX1 U9329 ( .A(n30635), .Y(n21067) );
  INVX1 U9330 ( .A(n29507), .Y(n21068) );
  INVX1 U9331 ( .A(n30073), .Y(n27019) );
  BUFX2 U9332 ( .A(n31901), .Y(n29209) );
  INVX1 U9333 ( .A(n26445), .Y(n26148) );
  INVX1 U9334 ( .A(n21023), .Y(n21069) );
  AND2X1 U9335 ( .A(n25779), .B(net89806), .Y(n30474) );
  AND2X2 U9336 ( .A(n30917), .B(net96340), .Y(n30928) );
  INVX1 U9337 ( .A(net112188), .Y(net150787) );
  BUFX2 U9338 ( .A(n3152), .Y(n21070) );
  INVX1 U9339 ( .A(n13804), .Y(n21071) );
  INVX1 U9340 ( .A(n30079), .Y(n21072) );
  INVX2 U9341 ( .A(n28597), .Y(n21097) );
  INVX1 U9342 ( .A(n29464), .Y(n21073) );
  INVX4 U9343 ( .A(n21095), .Y(n29464) );
  AND2X2 U9344 ( .A(n22994), .B(n22980), .Y(n21074) );
  INVX1 U9345 ( .A(n23091), .Y(n21076) );
  INVX1 U9346 ( .A(n21068), .Y(n23465) );
  MUX2X1 U9347 ( .B(n28388), .A(n28403), .S(n21077), .Y(n28406) );
  INVX1 U9348 ( .A(n26278), .Y(n21078) );
  INVX2 U9349 ( .A(n31894), .Y(n26278) );
  MUX2X1 U9350 ( .B(n28328), .A(n28327), .S(n21079), .Y(n28326) );
  MUX2X1 U9351 ( .B(n28475), .A(n28474), .S(n26514), .Y(n28473) );
  INVX1 U9352 ( .A(n26279), .Y(n21080) );
  INVX2 U9353 ( .A(n26446), .Y(n26096) );
  INVX2 U9354 ( .A(n26446), .Y(n26116) );
  INVX2 U9355 ( .A(n26446), .Y(n26115) );
  INVX2 U9356 ( .A(n26446), .Y(n26102) );
  INVX2 U9357 ( .A(n26446), .Y(n26127) );
  BUFX2 U9358 ( .A(grid[360]), .Y(n21081) );
  BUFX2 U9359 ( .A(grid[90]), .Y(n21082) );
  BUFX2 U9360 ( .A(grid[30]), .Y(n21083) );
  BUFX2 U9361 ( .A(grid[144]), .Y(n21084) );
  INVX1 U9362 ( .A(grid[6]), .Y(n21085) );
  INVX1 U9363 ( .A(n21085), .Y(n21086) );
  BUFX2 U9364 ( .A(grid[36]), .Y(n21087) );
  BUFX2 U9365 ( .A(grid[228]), .Y(n21088) );
  MUX2X1 U9366 ( .B(grid[210]), .A(grid[204]), .S(n26260), .Y(n28636) );
  INVX1 U9367 ( .A(n26113), .Y(n21089) );
  INVX2 U9368 ( .A(n26445), .Y(n26090) );
  MUX2X1 U9369 ( .B(n28514), .A(n28513), .S(n29461), .Y(n28512) );
  INVX4 U9370 ( .A(n29461), .Y(n28606) );
  INVX1 U9371 ( .A(n28596), .Y(n21090) );
  INVX1 U9372 ( .A(n28596), .Y(n21091) );
  INVX1 U9373 ( .A(n28596), .Y(n26516) );
  INVX1 U9374 ( .A(n31908), .Y(n21092) );
  INVX4 U9375 ( .A(alt5_net95668), .Y(net150650) );
  INVX4 U9376 ( .A(n29506), .Y(n25663) );
  BUFX2 U9377 ( .A(n25846), .Y(n21093) );
  AND2X2 U9378 ( .A(n23995), .B(n22022), .Y(n21818) );
  INVX1 U9379 ( .A(n21818), .Y(n21310) );
  MUX2X1 U9380 ( .B(n28556), .A(n28553), .S(n26304), .Y(n28560) );
  MUX2X1 U9381 ( .B(n28458), .A(n28457), .S(n21095), .Y(n28456) );
  INVX2 U9382 ( .A(n26162), .Y(n28597) );
  OAI21X1 U9383 ( .A(n29271), .B(n23382), .C(n21080), .Y(n21094) );
  INVX1 U9384 ( .A(n21094), .Y(n31500) );
  INVX4 U9385 ( .A(n8051), .Y(n21095) );
  INVX1 U9386 ( .A(n28595), .Y(n26121) );
  INVX2 U9387 ( .A(n28597), .Y(n26484) );
  INVX1 U9388 ( .A(n21095), .Y(n21096) );
  MUX2X1 U9389 ( .B(n28515), .A(n28518), .S(n21066), .Y(n28529) );
  NOR3X1 U9390 ( .A(n21099), .B(n32590), .C(n23464), .Y(n21098) );
  INVX2 U9391 ( .A(n21098), .Y(n32597) );
  INVX2 U9392 ( .A(n32591), .Y(n21099) );
  INVX1 U9393 ( .A(n29489), .Y(n21100) );
  INVX1 U9394 ( .A(n21100), .Y(n21101) );
  INVX1 U9395 ( .A(n21127), .Y(n33171) );
  INVX4 U9396 ( .A(n21103), .Y(n26445) );
  INVX4 U9397 ( .A(n25665), .Y(n28595) );
  MUX2X1 U9398 ( .B(n28561), .A(n28560), .S(n29461), .Y(n28559) );
  MUX2X1 U9399 ( .B(n25764), .A(n22688), .S(alt5_net95670), .Y(n8050) );
  INVX1 U9400 ( .A(alt5_net95668), .Y(alt5_net95662) );
  INVX1 U9401 ( .A(n8050), .Y(n21102) );
  INVX1 U9402 ( .A(n21102), .Y(n21103) );
  BUFX2 U9403 ( .A(n3772), .Y(n21104) );
  BUFX2 U9404 ( .A(n25668), .Y(n21105) );
  INVX2 U9405 ( .A(n34321), .Y(n34308) );
  OAI21X1 U9406 ( .A(n21108), .B(n25861), .C(n21109), .Y(n21107) );
  INVX1 U9407 ( .A(n34419), .Y(n21109) );
  INVX1 U9408 ( .A(n25861), .Y(n25862) );
  XOR2X1 U9409 ( .A(n21226), .B(n27913), .Y(n34386) );
  NOR3X1 U9410 ( .A(n34338), .B(n21111), .C(n34436), .Y(n21110) );
  INVX1 U9411 ( .A(n21110), .Y(n34438) );
  INVX1 U9412 ( .A(pLoc[2]), .Y(net110926) );
  INVX2 U9413 ( .A(net137490), .Y(alt14_net96238) );
  MUX2X1 U9414 ( .B(n25762), .A(n34248), .S(n23187), .Y(n21112) );
  BUFX2 U9415 ( .A(net110685), .Y(net150385) );
  INVX1 U9416 ( .A(net147983), .Y(net150376) );
  INVX4 U9417 ( .A(n29383), .Y(n29376) );
  INVX4 U9418 ( .A(n29383), .Y(n25466) );
  INVX1 U9419 ( .A(n26057), .Y(n21113) );
  INVX1 U9420 ( .A(net114253), .Y(net150330) );
  INVX1 U9421 ( .A(net150330), .Y(net150331) );
  INVX4 U9422 ( .A(n21209), .Y(n33682) );
  INVX2 U9423 ( .A(net105786), .Y(net110825) );
  INVX1 U9424 ( .A(net116949), .Y(net150253) );
  INVX1 U9425 ( .A(net105813), .Y(net116949) );
  INVX1 U9426 ( .A(alt14_net96264), .Y(net150251) );
  MUX2X1 U9427 ( .B(n28164), .A(n28165), .S(net105819), .Y(n28163) );
  INVX1 U9428 ( .A(n25645), .Y(n21114) );
  INVX1 U9429 ( .A(net150251), .Y(net150220) );
  MUX2X1 U9430 ( .B(n27984), .A(n27987), .S(net114744), .Y(n27991) );
  MUX2X1 U9431 ( .B(n28162), .A(n28161), .S(net149877), .Y(n28160) );
  INVX1 U9432 ( .A(oc[30]), .Y(n21115) );
  INVX4 U9433 ( .A(n21115), .Y(n21116) );
  MUX2X1 U9434 ( .B(grid[64]), .A(grid[70]), .S(net150132), .Y(n28210) );
  INVX4 U9435 ( .A(net109766), .Y(net150132) );
  INVX1 U9436 ( .A(n29602), .Y(n21117) );
  INVX1 U9437 ( .A(locTrig[1]), .Y(n29602) );
  INVX8 U9438 ( .A(net137490), .Y(net111222) );
  INVX4 U9439 ( .A(net150132), .Y(net150133) );
  MUX2X1 U9440 ( .B(grid[79]), .A(grid[73]), .S(net105857), .Y(n28024) );
  INVX1 U9441 ( .A(net150085), .Y(net150130) );
  INVX2 U9442 ( .A(net137490), .Y(net149947) );
  INVX1 U9443 ( .A(net150787), .Y(net150126) );
  INVX2 U9444 ( .A(net149909), .Y(net105857) );
  INVX1 U9445 ( .A(n21187), .Y(n15188) );
  INVX1 U9446 ( .A(alt14_net96248), .Y(net150085) );
  INVX1 U9447 ( .A(net149876), .Y(net105800) );
  INVX1 U9448 ( .A(net114244), .Y(net150046) );
  INVX1 U9449 ( .A(n29604), .Y(n21118) );
  AND2X2 U9450 ( .A(n22046), .B(n23925), .Y(n21843) );
  AND2X2 U9451 ( .A(n22050), .B(n23929), .Y(n21836) );
  INVX1 U9452 ( .A(n21833), .Y(n21298) );
  AND2X2 U9453 ( .A(n24012), .B(n22020), .Y(n21833) );
  MUX2X1 U9454 ( .B(grid[139]), .A(grid[133]), .S(net150787), .Y(n28016) );
  OAI21X1 U9455 ( .A(n24974), .B(n26055), .C(n33170), .Y(n21119) );
  OAI21X1 U9456 ( .A(n24262), .B(n34400), .C(n21147), .Y(n21120) );
  INVX1 U9457 ( .A(n21120), .Y(n34413) );
  INVX4 U9458 ( .A(n34411), .Y(n34400) );
  INVX1 U9459 ( .A(net149982), .Y(net149983) );
  MUX2X1 U9460 ( .B(grid[43]), .A(grid[37]), .S(net149922), .Y(n28031) );
  INVX1 U9461 ( .A(n21230), .Y(n21122) );
  NOR3X1 U9462 ( .A(n33166), .B(n26055), .C(n21122), .Y(n21121) );
  INVX1 U9463 ( .A(n21121), .Y(n33168) );
  NOR3X1 U9464 ( .A(n25401), .B(n26055), .C(n21230), .Y(n21123) );
  INVX1 U9465 ( .A(n21123), .Y(n33169) );
  INVX4 U9466 ( .A(n34434), .Y(n26055) );
  XNOR2X1 U9467 ( .A(n34393), .B(n25321), .Y(n21124) );
  NOR3X1 U9468 ( .A(locTrig[2]), .B(n22880), .C(n34612), .Y(n21125) );
  INVX1 U9469 ( .A(net109385), .Y(net149940) );
  INVX1 U9470 ( .A(net109385), .Y(net149941) );
  MUX2X1 U9471 ( .B(grid[236]), .A(grid[230]), .S(net150133), .Y(n28063) );
  INVX1 U9472 ( .A(net115535), .Y(net116925) );
  NOR3X1 U9473 ( .A(n25831), .B(n21229), .C(n21153), .Y(n21126) );
  INVX1 U9474 ( .A(n27178), .Y(n33068) );
  NOR3X1 U9475 ( .A(n34338), .B(n21128), .C(n21119), .Y(n21127) );
  INVX1 U9476 ( .A(net116776), .Y(net149922) );
  MUX2X1 U9477 ( .B(n28016), .A(n28015), .S(net105822), .Y(n28014) );
  OR2X2 U9478 ( .A(nc[10]), .B(nc[9]), .Y(n29547) );
  OAI21X1 U9479 ( .A(n25663), .B(n34187), .C(n21562), .Y(n21129) );
  INVX1 U9480 ( .A(n28603), .Y(n28604) );
  INVX1 U9481 ( .A(n28602), .Y(n28605) );
  MUX2X1 U9482 ( .B(n28031), .A(n28030), .S(net147761), .Y(n28029) );
  INVX2 U9483 ( .A(net105810), .Y(net147761) );
  INVX1 U9484 ( .A(net115635), .Y(net149876) );
  INVX1 U9485 ( .A(net115635), .Y(alt14_net96328) );
  MUX2X1 U9486 ( .B(n28037), .A(n28036), .S(n21130), .Y(n28035) );
  MUX2X1 U9487 ( .B(n27998), .A(n27997), .S(net147761), .Y(n27996) );
  XOR2X1 U9488 ( .A(n33079), .B(n33156), .Y(n25700) );
  BUFX2 U9489 ( .A(alt14_net96296), .Y(net149862) );
  BUFX2 U9490 ( .A(alt14_net96296), .Y(net149863) );
  INVX1 U9491 ( .A(alt14_net96302), .Y(alt14_net96296) );
  MUX2X1 U9492 ( .B(n28170), .A(n28171), .S(net105807), .Y(n28169) );
  MUX2X1 U9493 ( .B(n21132), .A(n21133), .S(n33113), .Y(n21131) );
  XNOR2X1 U9494 ( .A(n25855), .B(n25845), .Y(n21132) );
  XOR2X1 U9495 ( .A(n33112), .B(n23093), .Y(n21133) );
  INVX8 U9496 ( .A(n34305), .Y(n25759) );
  INVX1 U9497 ( .A(net109485), .Y(net149842) );
  INVX1 U9498 ( .A(n25730), .Y(n33100) );
  INVX1 U9499 ( .A(n20972), .Y(n21134) );
  INVX1 U9500 ( .A(pLoc[1]), .Y(net149749) );
  INVX1 U9501 ( .A(pLoc[1]), .Y(net95303) );
  OR2X2 U9502 ( .A(net151710), .B(n24973), .Y(n21135) );
  INVX4 U9503 ( .A(n29383), .Y(n29378) );
  INVX2 U9504 ( .A(n26043), .Y(n25850) );
  INVX1 U9505 ( .A(n22673), .Y(n25772) );
  INVX2 U9506 ( .A(n25150), .Y(n33573) );
  AND2X2 U9507 ( .A(n24009), .B(n22017), .Y(n21842) );
  INVX4 U9508 ( .A(n29383), .Y(n29377) );
  INVX1 U9509 ( .A(oc[1]), .Y(n21136) );
  INVX1 U9510 ( .A(n21201), .Y(n32745) );
  INVX1 U9511 ( .A(n21159), .Y(n21137) );
  INVX1 U9512 ( .A(n33068), .Y(n21138) );
  XOR2X1 U9513 ( .A(n25729), .B(n20969), .Y(n34352) );
  BUFX2 U9514 ( .A(n27218), .Y(n21139) );
  BUFX2 U9515 ( .A(oc[28]), .Y(n21140) );
  BUFX4 U9516 ( .A(oc[27]), .Y(n21141) );
  INVX2 U9517 ( .A(n25351), .Y(n33494) );
  AND2X2 U9518 ( .A(n26782), .B(n29612), .Y(n29617) );
  OR2X1 U9519 ( .A(oc[26]), .B(oc[28]), .Y(n29605) );
  INVX1 U9520 ( .A(n21843), .Y(n21289) );
  OR2X2 U9521 ( .A(n21164), .B(n21165), .Y(n33930) );
  INVX1 U9522 ( .A(n33930), .Y(n21142) );
  INVX1 U9523 ( .A(n29581), .Y(n21143) );
  OR2X2 U9524 ( .A(n21199), .B(n21200), .Y(n33708) );
  INVX1 U9525 ( .A(n33708), .Y(n21144) );
  BUFX2 U9526 ( .A(n32730), .Y(n21145) );
  BUFX2 U9527 ( .A(n32728), .Y(n21146) );
  NOR3X1 U9528 ( .A(n21148), .B(n21149), .C(n21150), .Y(n21147) );
  INVX1 U9529 ( .A(n34408), .Y(n21149) );
  INVX1 U9530 ( .A(n34409), .Y(n21150) );
  INVX1 U9531 ( .A(n21211), .Y(n29978) );
  AND2X2 U9532 ( .A(n25714), .B(n34356), .Y(n33134) );
  BUFX2 U9533 ( .A(pLoc[0]), .Y(n21151) );
  AND2X2 U9534 ( .A(n23286), .B(n25724), .Y(n21152) );
  INVX1 U9535 ( .A(n33068), .Y(n21153) );
  INVX1 U9536 ( .A(n21153), .Y(n21154) );
  INVX1 U9537 ( .A(n30626), .Y(n21155) );
  AND2X2 U9538 ( .A(n22047), .B(n23926), .Y(n21841) );
  INVX1 U9539 ( .A(net107091), .Y(net147983) );
  AND2X2 U9540 ( .A(n11954), .B(net96558), .Y(n21200) );
  AND2X2 U9541 ( .A(n26515), .B(n28602), .Y(n27272) );
  INVX1 U9542 ( .A(n29366), .Y(n21166) );
  INVX2 U9543 ( .A(alt5_net95670), .Y(alt5_net95654) );
  INVX2 U9544 ( .A(n21156), .Y(n27296) );
  AND2X2 U9545 ( .A(n32783), .B(n3181), .Y(n21157) );
  OR2X2 U9546 ( .A(n21157), .B(n21158), .Y(n22924) );
  OR2X2 U9547 ( .A(n22926), .B(n22925), .Y(n21158) );
  AND2X2 U9548 ( .A(n26066), .B(n23475), .Y(n21159) );
  AND2X1 U9549 ( .A(n26163), .B(n21186), .Y(n21195) );
  BUFX4 U9550 ( .A(n29685), .Y(n26163) );
  INVX2 U9551 ( .A(n33151), .Y(n33153) );
  INVX1 U9552 ( .A(n21841), .Y(n21291) );
  INVX1 U9553 ( .A(n27315), .Y(n21175) );
  AND2X2 U9554 ( .A(n29925), .B(n27315), .Y(n27303) );
  AND2X1 U9555 ( .A(n21211), .B(n27315), .Y(n29979) );
  INVX1 U9556 ( .A(oc[3]), .Y(n29723) );
  AND2X2 U9557 ( .A(n22045), .B(n23924), .Y(n21844) );
  INVX1 U9558 ( .A(n33021), .Y(n21160) );
  INVX1 U9559 ( .A(n22676), .Y(n33050) );
  XOR2X1 U9560 ( .A(n23201), .B(n34355), .Y(n34357) );
  INVX1 U9561 ( .A(n29383), .Y(n21161) );
  AND2X2 U9562 ( .A(n21219), .B(net96340), .Y(n21162) );
  INVX4 U9563 ( .A(n28597), .Y(n21163) );
  AND2X2 U9564 ( .A(n23280), .B(n33927), .Y(n21164) );
  AND2X2 U9565 ( .A(n27309), .B(n29423), .Y(n21165) );
  AND2X1 U9566 ( .A(n29037), .B(n2255), .Y(n25471) );
  MUX2X1 U9567 ( .B(grid[19]), .A(grid[13]), .S(net105857), .Y(n28034) );
  INVX1 U9568 ( .A(net116776), .Y(net116777) );
  MUX2X1 U9569 ( .B(n28063), .A(n28062), .S(net147761), .Y(n28061) );
  INVX4 U9570 ( .A(n21167), .Y(n29366) );
  INVX1 U9571 ( .A(n29385), .Y(n21167) );
  INVX1 U9572 ( .A(n29385), .Y(n29372) );
  INVX1 U9573 ( .A(n21844), .Y(n21288) );
  INVX1 U9574 ( .A(n8050), .Y(n26162) );
  AND2X2 U9575 ( .A(n29595), .B(n25421), .Y(n21168) );
  INVX1 U9576 ( .A(n26480), .Y(n26483) );
  INVX1 U9577 ( .A(n29379), .Y(n29382) );
  INVX4 U9578 ( .A(n29207), .Y(n29595) );
  INVX1 U9579 ( .A(n25205), .Y(n21169) );
  INVX1 U9580 ( .A(n34349), .Y(n21171) );
  INVX1 U9581 ( .A(n24989), .Y(n21172) );
  INVX1 U9582 ( .A(n26162), .Y(n21173) );
  NOR3X1 U9583 ( .A(n26939), .B(n23107), .C(n21175), .Y(n21174) );
  INVX1 U9584 ( .A(n26939), .Y(n29925) );
  INVX1 U9585 ( .A(n25753), .Y(n25714) );
  INVX1 U9586 ( .A(n21840), .Y(n21292) );
  NOR3X1 U9587 ( .A(n24127), .B(n33026), .C(n33025), .Y(n21177) );
  INVX8 U9588 ( .A(n21375), .Y(n33852) );
  BUFX2 U9589 ( .A(n21212), .Y(n21178) );
  INVX1 U9590 ( .A(n32706), .Y(n21179) );
  BUFX2 U9591 ( .A(n33016), .Y(n21180) );
  BUFX2 U9592 ( .A(n3164), .Y(n21181) );
  INVX1 U9593 ( .A(n25624), .Y(n29423) );
  INVX1 U9594 ( .A(n26304), .Y(n21231) );
  INVX2 U9595 ( .A(net90054), .Y(net147481) );
  INVX1 U9596 ( .A(net147481), .Y(net147490) );
  INVX1 U9597 ( .A(net147481), .Y(net147492) );
  INVX1 U9598 ( .A(net147481), .Y(net147493) );
  INVX1 U9599 ( .A(net147481), .Y(net147494) );
  INVX1 U9600 ( .A(net147481), .Y(net147495) );
  INVX1 U9601 ( .A(net147493), .Y(net147496) );
  INVX1 U9602 ( .A(net147490), .Y(net147497) );
  INVX1 U9603 ( .A(net147493), .Y(net147498) );
  INVX1 U9604 ( .A(net147492), .Y(net147499) );
  INVX1 U9605 ( .A(net147494), .Y(net147500) );
  INVX1 U9606 ( .A(net147494), .Y(net147501) );
  INVX1 U9607 ( .A(net147495), .Y(net147502) );
  INVX1 U9608 ( .A(net151741), .Y(net147504) );
  INVX1 U9609 ( .A(net147492), .Y(net147505) );
  INVX1 U9610 ( .A(net147495), .Y(net147507) );
  INVX1 U9611 ( .A(net110814), .Y(net110815) );
  INVX2 U9612 ( .A(net110814), .Y(net147379) );
  INVX4 U9613 ( .A(n21185), .Y(n21186) );
  INVX1 U9614 ( .A(n21203), .Y(n21182) );
  INVX2 U9615 ( .A(n21182), .Y(n21183) );
  INVX1 U9616 ( .A(n21182), .Y(n21185) );
  MUX2X1 U9617 ( .B(n25326), .A(n25725), .S(n34252), .Y(n34238) );
  NOR3X1 U9618 ( .A(n21024), .B(n29489), .C(n21028), .Y(n21187) );
  AND2X1 U9619 ( .A(n32653), .B(n32652), .Y(n32654) );
  AND2X2 U9620 ( .A(n9141), .B(n29381), .Y(n21798) );
  INVX1 U9621 ( .A(n32738), .Y(n21202) );
  AND2X2 U9622 ( .A(n23299), .B(n25724), .Y(n21188) );
  INVX1 U9623 ( .A(net111205), .Y(net110814) );
  INVX1 U9624 ( .A(n26078), .Y(n26521) );
  NOR3X1 U9625 ( .A(n21190), .B(n32833), .C(n24793), .Y(n21189) );
  INVX1 U9626 ( .A(n21189), .Y(n32840) );
  INVX1 U9627 ( .A(n32832), .Y(n21190) );
  INVX1 U9628 ( .A(n25114), .Y(n21191) );
  INVX1 U9629 ( .A(alt5_net95668), .Y(net113321) );
  INVX1 U9630 ( .A(n27058), .Y(n21192) );
  AND2X2 U9631 ( .A(n30186), .B(n21193), .Y(n25715) );
  AND2X1 U9632 ( .A(n21195), .B(n30281), .Y(n21193) );
  INVX1 U9633 ( .A(n26050), .Y(n21194) );
  NOR3X1 U9634 ( .A(n21197), .B(n24442), .C(n20848), .Y(n21196) );
  INVX1 U9635 ( .A(n30049), .Y(n21197) );
  INVX1 U9636 ( .A(n25079), .Y(n21198) );
  AND2X2 U9637 ( .A(n29399), .B(n33718), .Y(n21199) );
  INVX1 U9638 ( .A(n26050), .Y(n29504) );
  INVX4 U9639 ( .A(n29401), .Y(n29399) );
  NOR3X1 U9640 ( .A(n24790), .B(n32737), .C(n21202), .Y(n21201) );
  XNOR2X1 U9641 ( .A(n25859), .B(n34442), .Y(n34233) );
  INVX2 U9642 ( .A(n26337), .Y(n26339) );
  INVX4 U9643 ( .A(n21173), .Y(n26446) );
  INVX1 U9644 ( .A(n21163), .Y(n26139) );
  INVX1 U9645 ( .A(loc_s2[3]), .Y(n21205) );
  INVX1 U9646 ( .A(n13706), .Y(n21206) );
  OAI21X1 U9647 ( .A(n21204), .B(n21205), .C(n21206), .Y(n21203) );
  INVX1 U9648 ( .A(n13799), .Y(n29626) );
  OAI21X1 U9649 ( .A(n21208), .B(n21204), .C(n13707), .Y(n21207) );
  NOR3X1 U9650 ( .A(n27081), .B(n21175), .C(n23108), .Y(n21209) );
  INVX4 U9651 ( .A(n23108), .Y(n29835) );
  NOR3X1 U9652 ( .A(locTrig[2]), .B(n22880), .C(n21170), .Y(n21210) );
  NOR3X1 U9653 ( .A(oc[2]), .B(oc[1]), .C(oc[0]), .Y(n21211) );
  INVX1 U9654 ( .A(oc[2]), .Y(n29745) );
  INVX1 U9655 ( .A(oc[1]), .Y(n29756) );
  AND2X1 U9656 ( .A(n22044), .B(n21514), .Y(n24886) );
  INVX1 U9657 ( .A(n26810), .Y(n21212) );
  INVX1 U9658 ( .A(n27912), .Y(n21227) );
  OAI21X1 U9659 ( .A(n29271), .B(n23396), .C(n26281), .Y(n21213) );
  INVX1 U9660 ( .A(n21213), .Y(n31636) );
  OAI21X1 U9661 ( .A(n29271), .B(n23420), .C(n26281), .Y(n21214) );
  INVX1 U9662 ( .A(n21214), .Y(n31849) );
  BUFX2 U9663 ( .A(grid[367]), .Y(n21215) );
  AND2X2 U9664 ( .A(n30186), .B(n21216), .Y(n25720) );
  AND2X1 U9665 ( .A(n30281), .B(n20977), .Y(n21216) );
  INVX1 U9666 ( .A(n26270), .Y(n21217) );
  OAI21X1 U9667 ( .A(n29271), .B(n23375), .C(n26277), .Y(n21218) );
  INVX1 U9668 ( .A(n21218), .Y(n31442) );
  AND2X2 U9669 ( .A(net109585), .B(net125066), .Y(n21219) );
  INVX1 U9670 ( .A(n26869), .Y(n21220) );
  INVX1 U9671 ( .A(n26869), .Y(n32877) );
  INVX2 U9672 ( .A(locTrig[3]), .Y(n29484) );
  MUX2X1 U9673 ( .B(n28503), .A(n28500), .S(n29462), .Y(n28514) );
  AND2X2 U9674 ( .A(n30033), .B(n3209), .Y(n21221) );
  OR2X2 U9675 ( .A(n26797), .B(n25634), .Y(n21222) );
  INVX4 U9676 ( .A(n26797), .Y(n30033) );
  MUX2X1 U9677 ( .B(n28366), .A(n28365), .S(n21095), .Y(n28364) );
  INVX1 U9678 ( .A(n28595), .Y(n26122) );
  INVX1 U9679 ( .A(oc[2]), .Y(n21223) );
  INVX4 U9680 ( .A(n21223), .Y(n21224) );
  AND2X2 U9681 ( .A(n24010), .B(n22018), .Y(n21838) );
  INVX1 U9682 ( .A(n21836), .Y(n21296) );
  OR2X2 U9683 ( .A(n32756), .B(n32755), .Y(n32763) );
  AND2X2 U9684 ( .A(n23944), .B(n22078), .Y(n21845) );
  INVX1 U9685 ( .A(n23091), .Y(n29507) );
  AND2X2 U9686 ( .A(n30281), .B(n26339), .Y(n27310) );
  BUFX2 U9687 ( .A(n34209), .Y(n25615) );
  INVX1 U9688 ( .A(n26270), .Y(n26272) );
  XNOR2X1 U9689 ( .A(n29475), .B(n2255), .Y(n21225) );
  INVX2 U9690 ( .A(n21225), .Y(n27318) );
  INVX1 U9691 ( .A(n2253), .Y(n26051) );
  INVX2 U9692 ( .A(n27904), .Y(n27907) );
  OR2X2 U9693 ( .A(n34380), .B(n21227), .Y(n21226) );
  AND2X2 U9694 ( .A(n24011), .B(n22019), .Y(n21837) );
  INVX1 U9695 ( .A(n29382), .Y(n29380) );
  AND2X2 U9696 ( .A(n22992), .B(n25849), .Y(n21228) );
  INVX4 U9697 ( .A(n27905), .Y(n27908) );
  INVX4 U9698 ( .A(alt5_net95670), .Y(alt5_net95658) );
  INVX4 U9699 ( .A(n22940), .Y(n33908) );
  INVX1 U9700 ( .A(n21837), .Y(n21295) );
  AND2X2 U9701 ( .A(oc[16]), .B(n27316), .Y(n29719) );
  INVX1 U9702 ( .A(n21426), .Y(n21229) );
  AND2X2 U9703 ( .A(n26045), .B(n23098), .Y(n21230) );
  INVX4 U9704 ( .A(n15188), .Y(n29506) );
  MUX2X1 U9705 ( .B(n28521), .A(n28524), .S(n29463), .Y(n28528) );
  MUX2X1 U9706 ( .B(n28487), .A(n28486), .S(n26514), .Y(n28485) );
  MUX2X1 U9707 ( .B(grid[58]), .A(grid[52]), .S(n21097), .Y(n28519) );
  MUX2X1 U9708 ( .B(n28526), .A(n28525), .S(n28599), .Y(n28524) );
  MUX2X1 U9709 ( .B(n25405), .A(n25664), .S(n25653), .Y(n34393) );
  AND2X2 U9710 ( .A(n32936), .B(n32935), .Y(n32937) );
  AND2X2 U9711 ( .A(n29719), .B(n23922), .Y(n29720) );
  AND2X2 U9712 ( .A(n26838), .B(n29604), .Y(n29609) );
  INVX1 U9713 ( .A(n21842), .Y(n21290) );
  AND2X2 U9714 ( .A(oc[14]), .B(oc[12]), .Y(n27316) );
  AND2X1 U9715 ( .A(n33326), .B(n3247), .Y(n32918) );
  INVX1 U9716 ( .A(n21831), .Y(n21300) );
  AND2X2 U9717 ( .A(n22057), .B(n23932), .Y(n21831) );
  AND2X2 U9718 ( .A(n22070), .B(n23938), .Y(n21824) );
  INVX4 U9719 ( .A(n33682), .Y(n33696) );
  AND2X2 U9720 ( .A(n23288), .B(n30626), .Y(n21232) );
  INVX1 U9721 ( .A(n34373), .Y(n21233) );
  NOR3X1 U9722 ( .A(n24124), .B(n32729), .C(n21235), .Y(n21234) );
  INVX1 U9723 ( .A(n21234), .Y(n32735) );
  INVX1 U9724 ( .A(net112858), .Y(net146838) );
  AND2X2 U9725 ( .A(n25688), .B(n20974), .Y(n21236) );
  OR2X2 U9726 ( .A(net151977), .B(n21238), .Y(n21237) );
  OR2X2 U9727 ( .A(n22963), .B(n21237), .Y(net146826) );
  INVX1 U9728 ( .A(n21838), .Y(n21294) );
  INVX1 U9729 ( .A(n21825), .Y(n21306) );
  AND2X2 U9730 ( .A(net144199), .B(n23937), .Y(n21825) );
  INVX1 U9731 ( .A(n21827), .Y(n21304) );
  AND2X2 U9732 ( .A(n23935), .B(n22065), .Y(n21827) );
  INVX4 U9733 ( .A(n25753), .Y(n25688) );
  INVX1 U9734 ( .A(n21845), .Y(n21311) );
  INVX1 U9735 ( .A(n21824), .Y(n21307) );
  INVX1 U9736 ( .A(n21322), .Y(n21239) );
  OR2X2 U9737 ( .A(n22094), .B(n25479), .Y(n11049) );
  AND2X2 U9738 ( .A(n23949), .B(n21995), .Y(n21318) );
  INVX1 U9739 ( .A(n21318), .Y(n21242) );
  AND2X2 U9740 ( .A(n23951), .B(n20976), .Y(n21317) );
  INVX1 U9741 ( .A(n21317), .Y(n21243) );
  AND2X2 U9742 ( .A(n23953), .B(n23898), .Y(n21316) );
  INVX1 U9743 ( .A(n21316), .Y(n21244) );
  AND2X2 U9744 ( .A(n23955), .B(n23900), .Y(n21315) );
  INVX1 U9745 ( .A(n21315), .Y(n21245) );
  AND2X2 U9746 ( .A(n23957), .B(n23901), .Y(n21314) );
  INVX1 U9747 ( .A(n21314), .Y(n21246) );
  OR2X2 U9748 ( .A(n25345), .B(n33175), .Y(n21860) );
  INVX1 U9749 ( .A(n21860), .Y(n21247) );
  AND2X2 U9750 ( .A(n23960), .B(n21996), .Y(n21521) );
  INVX1 U9751 ( .A(n21521), .Y(n21248) );
  AND2X2 U9752 ( .A(n23961), .B(n22026), .Y(n21513) );
  INVX1 U9753 ( .A(n21513), .Y(n21249) );
  AND2X2 U9754 ( .A(n23962), .B(n33452), .Y(n21512) );
  INVX1 U9755 ( .A(n21512), .Y(n21250) );
  AND2X2 U9756 ( .A(n23963), .B(n33469), .Y(n21504) );
  INVX1 U9757 ( .A(n21504), .Y(n21251) );
  AND2X2 U9758 ( .A(n23964), .B(n33475), .Y(n21503) );
  INVX1 U9759 ( .A(n21503), .Y(n21252) );
  AND2X2 U9760 ( .A(n22027), .B(n23965), .Y(n21495) );
  INVX1 U9761 ( .A(n21495), .Y(n21253) );
  AND2X2 U9762 ( .A(n23966), .B(n22028), .Y(n21494) );
  INVX1 U9763 ( .A(n21494), .Y(n21254) );
  AND2X2 U9764 ( .A(n23967), .B(n22029), .Y(n21486) );
  INVX1 U9765 ( .A(n21486), .Y(n21255) );
  AND2X2 U9766 ( .A(n23968), .B(n33521), .Y(n21485) );
  INVX1 U9767 ( .A(n21485), .Y(n21256) );
  AND2X2 U9768 ( .A(n23969), .B(n22030), .Y(n21468) );
  INVX1 U9769 ( .A(n21468), .Y(n21257) );
  AND2X2 U9770 ( .A(n22031), .B(n23970), .Y(n21466) );
  INVX1 U9771 ( .A(n21466), .Y(n21258) );
  AND2X2 U9772 ( .A(n23971), .B(n22032), .Y(n21458) );
  INVX1 U9773 ( .A(n21458), .Y(n21259) );
  AND2X2 U9774 ( .A(n23972), .B(n22033), .Y(n21457) );
  INVX1 U9775 ( .A(n21457), .Y(n21260) );
  AND2X2 U9776 ( .A(n23973), .B(n33616), .Y(n21449) );
  INVX1 U9777 ( .A(n21449), .Y(n21261) );
  AND2X2 U9778 ( .A(n23974), .B(n22034), .Y(n21448) );
  INVX1 U9779 ( .A(n21448), .Y(n21262) );
  AND2X2 U9780 ( .A(n23975), .B(n22035), .Y(n21440) );
  INVX1 U9781 ( .A(n21440), .Y(n21263) );
  AND2X2 U9782 ( .A(n23976), .B(n22036), .Y(n21439) );
  INVX1 U9783 ( .A(n21439), .Y(n21264) );
  AND2X2 U9784 ( .A(n23977), .B(n22037), .Y(n21431) );
  INVX1 U9785 ( .A(n21431), .Y(n21265) );
  AND2X2 U9786 ( .A(n23978), .B(n22038), .Y(n21430) );
  INVX1 U9787 ( .A(n21430), .Y(n21266) );
  AND2X2 U9788 ( .A(n23979), .B(n21997), .Y(n21422) );
  INVX1 U9789 ( .A(n21422), .Y(n21267) );
  AND2X2 U9790 ( .A(n23980), .B(n21998), .Y(n21421) );
  INVX1 U9791 ( .A(n21421), .Y(n21268) );
  AND2X2 U9792 ( .A(n23999), .B(n21999), .Y(n21413) );
  INVX1 U9793 ( .A(n21413), .Y(n21269) );
  AND2X2 U9794 ( .A(n21144), .B(n23981), .Y(n21412) );
  INVX1 U9795 ( .A(n21412), .Y(n21270) );
  AND2X2 U9796 ( .A(n23982), .B(n22000), .Y(n21404) );
  AND2X2 U9797 ( .A(n22001), .B(n23983), .Y(n21403) );
  INVX1 U9798 ( .A(n21403), .Y(n21272) );
  AND2X2 U9799 ( .A(n23984), .B(n22002), .Y(n21395) );
  INVX1 U9800 ( .A(n21395), .Y(n21273) );
  AND2X2 U9801 ( .A(n24000), .B(n22003), .Y(n21394) );
  INVX1 U9802 ( .A(n21394), .Y(n21274) );
  AND2X2 U9803 ( .A(n23985), .B(n22004), .Y(n21386) );
  INVX1 U9804 ( .A(n21386), .Y(n21275) );
  AND2X2 U9805 ( .A(n23986), .B(n22005), .Y(n21385) );
  INVX1 U9806 ( .A(n21385), .Y(n21276) );
  AND2X2 U9807 ( .A(n23987), .B(n22006), .Y(n21377) );
  INVX1 U9808 ( .A(n21377), .Y(n21277) );
  AND2X2 U9809 ( .A(n23988), .B(n22007), .Y(n21376) );
  INVX1 U9810 ( .A(n21376), .Y(n21278) );
  AND2X2 U9811 ( .A(n24001), .B(n22008), .Y(n21368) );
  INVX1 U9812 ( .A(n21368), .Y(n21279) );
  AND2X2 U9813 ( .A(n24002), .B(n22009), .Y(n21367) );
  INVX1 U9814 ( .A(n21367), .Y(n21280) );
  AND2X2 U9815 ( .A(n23989), .B(n22010), .Y(n21359) );
  INVX1 U9816 ( .A(n21359), .Y(n21281) );
  AND2X2 U9817 ( .A(n23990), .B(n22011), .Y(n21358) );
  INVX1 U9818 ( .A(n21358), .Y(n21282) );
  AND2X2 U9819 ( .A(n23991), .B(n22012), .Y(n21350) );
  INVX1 U9820 ( .A(n21350), .Y(n21283) );
  AND2X2 U9821 ( .A(n23992), .B(n22013), .Y(n21349) );
  INVX1 U9822 ( .A(n21349), .Y(n21284) );
  AND2X2 U9823 ( .A(n23993), .B(n22014), .Y(n21341) );
  INVX1 U9824 ( .A(n21341), .Y(n21285) );
  AND2X2 U9825 ( .A(n24003), .B(n22015), .Y(n21340) );
  INVX1 U9826 ( .A(n21340), .Y(n21286) );
  AND2X2 U9827 ( .A(n23994), .B(n22016), .Y(n20535) );
  INVX1 U9828 ( .A(n20535), .Y(n21287) );
  AND2X1 U9829 ( .A(n22049), .B(n23928), .Y(n21839) );
  AND2X2 U9830 ( .A(n22051), .B(n23930), .Y(n21835) );
  INVX1 U9831 ( .A(n21835), .Y(n21297) );
  AND2X2 U9832 ( .A(n22061), .B(n23933), .Y(n21830) );
  INVX1 U9833 ( .A(n21830), .Y(n21301) );
  AND2X1 U9834 ( .A(n22062), .B(n23934), .Y(n21829) );
  AND2X2 U9835 ( .A(n24013), .B(n22021), .Y(n21828) );
  INVX1 U9836 ( .A(n21828), .Y(n21303) );
  AND2X1 U9837 ( .A(n22069), .B(n23936), .Y(n21826) );
  AND2X1 U9838 ( .A(n22073), .B(n23941), .Y(n21821) );
  AND2X2 U9839 ( .A(n22077), .B(n23942), .Y(n21819) );
  INVX1 U9840 ( .A(n21819), .Y(n21309) );
  AND2X2 U9841 ( .A(n23996), .B(n22023), .Y(n21816) );
  INVX1 U9842 ( .A(n21816), .Y(n21312) );
  OR2X2 U9843 ( .A(n33995), .B(n29363), .Y(n21603) );
  INVX1 U9844 ( .A(n21603), .Y(n21319) );
  OR2X1 U9845 ( .A(n29370), .B(n34029), .Y(n21637) );
  INVX1 U9846 ( .A(n21637), .Y(n21320) );
  OR2X1 U9847 ( .A(n29370), .B(n34042), .Y(n21650) );
  INVX1 U9848 ( .A(n21650), .Y(n21321) );
  OR2X1 U9849 ( .A(n29365), .B(n34055), .Y(n21663) );
  INVX1 U9850 ( .A(n21663), .Y(n21326) );
  OR2X1 U9851 ( .A(n29370), .B(n34068), .Y(n21677) );
  INVX1 U9852 ( .A(n21677), .Y(n21327) );
  OR2X1 U9853 ( .A(n29371), .B(n34081), .Y(n21690) );
  INVX1 U9854 ( .A(n21690), .Y(n21330) );
  OR2X1 U9855 ( .A(n29371), .B(n34094), .Y(n21704) );
  INVX1 U9856 ( .A(n21704), .Y(n21333) );
  OR2X1 U9857 ( .A(n29366), .B(n34107), .Y(n21717) );
  INVX1 U9858 ( .A(n21717), .Y(n21336) );
  OR2X1 U9859 ( .A(n29367), .B(n34120), .Y(n21730) );
  INVX1 U9860 ( .A(n21730), .Y(n21339) );
  OR2X1 U9861 ( .A(n29368), .B(n34133), .Y(n21743) );
  INVX1 U9862 ( .A(n21743), .Y(n21342) );
  OR2X2 U9863 ( .A(n29369), .B(n34146), .Y(n21756) );
  INVX1 U9864 ( .A(n21756), .Y(n21345) );
  AND2X2 U9865 ( .A(n22081), .B(n23902), .Y(n20538) );
  INVX1 U9866 ( .A(n20538), .Y(n21348) );
  AND2X2 U9867 ( .A(n23997), .B(n22024), .Y(n20536) );
  INVX1 U9868 ( .A(n20536), .Y(n21351) );
  OR2X2 U9869 ( .A(n34231), .B(n25345), .Y(n21854) );
  INVX1 U9870 ( .A(n30638), .Y(n30079) );
  OR2X2 U9871 ( .A(n25590), .B(n23347), .Y(n25591) );
  INVX1 U9872 ( .A(n25591), .Y(n21357) );
  OR2X2 U9873 ( .A(n32470), .B(n32469), .Y(n25747) );
  INVX1 U9874 ( .A(n25747), .Y(n21360) );
  AND2X2 U9875 ( .A(n25839), .B(n34385), .Y(n25835) );
  INVX1 U9876 ( .A(n25835), .Y(n21363) );
  OR2X2 U9877 ( .A(nc[1]), .B(n22142), .Y(n29552) );
  INVX1 U9878 ( .A(n29552), .Y(n21366) );
  OR2X2 U9879 ( .A(n27196), .B(n33928), .Y(n29566) );
  INVX1 U9880 ( .A(n29566), .Y(n21369) );
  INVX1 U9881 ( .A(n29979), .Y(n21372) );
  AND2X2 U9882 ( .A(n29835), .B(n23445), .Y(n33837) );
  AND2X2 U9883 ( .A(n29835), .B(n23297), .Y(n33770) );
  AND2X2 U9884 ( .A(n29831), .B(n27315), .Y(n30024) );
  INVX1 U9885 ( .A(n30024), .Y(n21381) );
  AND2X2 U9886 ( .A(n30626), .B(n23283), .Y(n33398) );
  AND2X2 U9887 ( .A(n30626), .B(n29902), .Y(n33215) );
  AND2X2 U9888 ( .A(n23448), .B(n29330), .Y(n32479) );
  INVX1 U9889 ( .A(n32479), .Y(n21390) );
  AND2X2 U9890 ( .A(n25878), .B(n32387), .Y(n31528) );
  INVX1 U9891 ( .A(n31528), .Y(n21393) );
  OR2X2 U9892 ( .A(n21155), .B(n32970), .Y(n32972) );
  INVX1 U9893 ( .A(n32972), .Y(n21396) );
  OR2X1 U9894 ( .A(n27911), .B(n25864), .Y(n34376) );
  INVX1 U9895 ( .A(n34376), .Y(n21399) );
  OR2X2 U9896 ( .A(n20812), .B(n27192), .Y(n14674) );
  INVX1 U9897 ( .A(n14674), .Y(n21402) );
  OR2X2 U9898 ( .A(n22885), .B(n22886), .Y(n22883) );
  OR2X2 U9899 ( .A(n22884), .B(n32503), .Y(n22886) );
  OR2X2 U9900 ( .A(n22891), .B(n22892), .Y(n22889) );
  OR2X2 U9901 ( .A(n22890), .B(n32579), .Y(n22892) );
  OR2X2 U9902 ( .A(n22894), .B(n22895), .Y(n22893) );
  OR2X2 U9903 ( .A(n24782), .B(n32599), .Y(n22895) );
  OR2X2 U9904 ( .A(n22899), .B(n22900), .Y(n22897) );
  OR2X2 U9905 ( .A(n22898), .B(n32682), .Y(n22900) );
  OR2X2 U9906 ( .A(n22903), .B(n22904), .Y(n22901) );
  OR2X2 U9907 ( .A(n32691), .B(n22902), .Y(n22904) );
  OR2X2 U9908 ( .A(n22909), .B(n32788), .Y(n22906) );
  OR2X2 U9909 ( .A(n22907), .B(n22908), .Y(n22909) );
  OR2X2 U9910 ( .A(n22912), .B(n22913), .Y(n22910) );
  OR2X2 U9911 ( .A(n22911), .B(n32860), .Y(n22913) );
  OR2X2 U9912 ( .A(n22916), .B(n22917), .Y(n22914) );
  OR2X2 U9913 ( .A(n22915), .B(n32868), .Y(n22917) );
  OR2X2 U9914 ( .A(n22922), .B(n22923), .Y(n22920) );
  OR2X2 U9915 ( .A(n22921), .B(n32959), .Y(n22923) );
  OR2X2 U9916 ( .A(n22936), .B(n22937), .Y(n22934) );
  OR2X2 U9917 ( .A(n22935), .B(n32779), .Y(n22937) );
  OR2X2 U9918 ( .A(net143109), .B(net138174), .Y(n22963) );
  OR2X2 U9919 ( .A(n22977), .B(n22978), .Y(n22975) );
  OR2X2 U9920 ( .A(n22976), .B(n32879), .Y(n22978) );
  OR2X2 U9921 ( .A(n23212), .B(n21016), .Y(n23211) );
  OR2X2 U9922 ( .A(n23215), .B(n21021), .Y(n23214) );
  OR2X2 U9923 ( .A(n23218), .B(n21025), .Y(n23217) );
  OR2X2 U9924 ( .A(n23225), .B(n23226), .Y(n23223) );
  OR2X2 U9925 ( .A(n23224), .B(n30759), .Y(n23226) );
  OR2X2 U9926 ( .A(n23228), .B(n21036), .Y(n23227) );
  OR2X2 U9927 ( .A(n23232), .B(n23233), .Y(n23230) );
  OR2X2 U9928 ( .A(n23231), .B(n30799), .Y(n23233) );
  OR2X2 U9929 ( .A(n23238), .B(n21017), .Y(n23237) );
  OR2X2 U9930 ( .A(n23241), .B(n21034), .Y(n23240) );
  OR2X2 U9931 ( .A(n23244), .B(n20830), .Y(n23243) );
  OR2X2 U9932 ( .A(n23247), .B(n21035), .Y(n23246) );
  OR2X2 U9933 ( .A(n23250), .B(n21026), .Y(n23249) );
  OR2X2 U9934 ( .A(n23253), .B(n21010), .Y(n23252) );
  OR2X2 U9935 ( .A(n23257), .B(n23258), .Y(n23255) );
  OR2X2 U9936 ( .A(n23256), .B(n31543), .Y(n23258) );
  OR2X2 U9937 ( .A(n23260), .B(n21014), .Y(n23259) );
  OR2X2 U9938 ( .A(n23264), .B(n23265), .Y(n23262) );
  OR2X2 U9939 ( .A(n23263), .B(n31678), .Y(n23265) );
  OR2X2 U9940 ( .A(n23267), .B(n21015), .Y(n23266) );
  OR2X2 U9941 ( .A(n23271), .B(n23272), .Y(n23269) );
  OR2X2 U9942 ( .A(n24711), .B(n23270), .Y(n23272) );
  OR2X2 U9943 ( .A(n23618), .B(n20835), .Y(n23617) );
  OR2X2 U9944 ( .A(n23621), .B(n21018), .Y(n23620) );
  OR2X2 U9945 ( .A(n23624), .B(n21019), .Y(n23623) );
  OR2X2 U9946 ( .A(n23637), .B(n23638), .Y(n23634) );
  INVX1 U9947 ( .A(n23634), .Y(n21405) );
  OR2X2 U9948 ( .A(n23635), .B(n23636), .Y(n23638) );
  AND2X2 U9949 ( .A(n23437), .B(n23435), .Y(n24880) );
  AND2X2 U9950 ( .A(n23959), .B(n23923), .Y(n24881) );
  AND2X2 U9951 ( .A(n22042), .B(n21508), .Y(n24884) );
  AND2X2 U9952 ( .A(n22043), .B(n22040), .Y(n24885) );
  AND2X1 U9953 ( .A(n27223), .B(net96340), .Y(n24936) );
  AND2X2 U9954 ( .A(n34385), .B(n26978), .Y(n24984) );
  INVX1 U9955 ( .A(n24984), .Y(n21411) );
  OR2X2 U9956 ( .A(n26339), .B(n24991), .Y(n24989) );
  INVX1 U9957 ( .A(n24989), .Y(n21414) );
  OR2X2 U9958 ( .A(n24990), .B(n21186), .Y(n24991) );
  AND2X2 U9959 ( .A(T[1]), .B(n34375), .Y(n25195) );
  OR2X2 U9960 ( .A(n25318), .B(n25319), .Y(n25320) );
  OR2X2 U9961 ( .A(n25460), .B(n31513), .Y(n25461) );
  AND2X2 U9962 ( .A(n24005), .B(n24006), .Y(n25472) );
  OR2X2 U9963 ( .A(n31783), .B(n29277), .Y(n25477) );
  OR2X2 U9964 ( .A(n22097), .B(n25477), .Y(n31780) );
  INVX1 U9965 ( .A(n31780), .Y(n21417) );
  OR2X1 U9966 ( .A(n34340), .B(n34338), .Y(n25479) );
  OR2X2 U9967 ( .A(n32822), .B(n32821), .Y(n25517) );
  AND2X2 U9968 ( .A(n24007), .B(n23603), .Y(n25524) );
  AND2X2 U9969 ( .A(n24008), .B(n23918), .Y(n25527) );
  OR2X2 U9970 ( .A(n27064), .B(n23207), .Y(n29600) );
  AND2X2 U9971 ( .A(n25569), .B(n25570), .Y(n25571) );
  INVX1 U9972 ( .A(n25571), .Y(n21420) );
  OR2X2 U9973 ( .A(n31650), .B(n31648), .Y(n25606) );
  OR2X1 U9974 ( .A(n25754), .B(n34338), .Y(n25662) );
  OR2X2 U9975 ( .A(n25728), .B(T[0]), .Y(n25664) );
  OR2X2 U9976 ( .A(n31614), .B(n31612), .Y(n25669) );
  OR2X2 U9977 ( .A(n25859), .B(T[3]), .Y(n25725) );
  AND2X2 U9978 ( .A(T[4]), .B(n33077), .Y(n25726) );
  OR2X2 U9979 ( .A(n13800), .B(n29626), .Y(n25778) );
  OR2X2 U9980 ( .A(n34357), .B(n34356), .Y(n25849) );
  OR2X2 U9981 ( .A(n33062), .B(T[0]), .Y(n25855) );
  AND2X2 U9982 ( .A(n29619), .B(n29618), .Y(n26066) );
  AND2X2 U9983 ( .A(n22086), .B(n23920), .Y(n27042) );
  AND2X2 U9984 ( .A(n3161), .B(n23450), .Y(n27142) );
  INVX1 U9985 ( .A(n27142), .Y(n21423) );
  OR2X2 U9986 ( .A(n23080), .B(n25575), .Y(n29189) );
  INVX1 U9987 ( .A(n29189), .Y(n21426) );
  AND2X2 U9988 ( .A(n29603), .B(n21134), .Y(net90053) );
  AND2X2 U9989 ( .A(Setup[0]), .B(net90053), .Y(n16281) );
  AND2X2 U9990 ( .A(n23074), .B(n24978), .Y(net53176) );
  AND2X2 U9991 ( .A(n2255), .B(n2254), .Y(n29479) );
  AND2X2 U9992 ( .A(n23200), .B(n25335), .Y(n29575) );
  AND2X2 U9993 ( .A(n27196), .B(n23200), .Y(n29590) );
  AND2X2 U9994 ( .A(n22041), .B(n21994), .Y(n13708) );
  AND2X2 U9995 ( .A(n21172), .B(n30410), .Y(n32042) );
  INVX1 U9996 ( .A(net95147), .Y(net145105) );
  AND2X2 U9997 ( .A(n23946), .B(n29631), .Y(n30486) );
  INVX1 U9998 ( .A(n30486), .Y(n21429) );
  AND2X2 U9999 ( .A(Setup[1]), .B(n16281), .Y(n30656) );
  AND2X2 U10000 ( .A(net90053), .B(n29704), .Y(n30657) );
  INVX1 U10001 ( .A(n30657), .Y(n21432) );
  AND2X2 U10002 ( .A(n23285), .B(n30626), .Y(n33638) );
  AND2X2 U10003 ( .A(n23290), .B(n30626), .Y(n33595) );
  AND2X2 U10004 ( .A(n29993), .B(n21106), .Y(n33019) );
  AND2X2 U10005 ( .A(n23291), .B(n29331), .Y(n32783) );
  AND2X2 U10006 ( .A(n23293), .B(n30626), .Y(n33572) );
  AND2X2 U10007 ( .A(n23295), .B(n30626), .Y(n32553) );
  AND2X2 U10008 ( .A(n29807), .B(n30626), .Y(n33493) );
  AND2X2 U10009 ( .A(n30040), .B(n21106), .Y(n32528) );
  AND2X2 U10010 ( .A(n23299), .B(n30626), .Y(n33470) );
  AND2X2 U10011 ( .A(n23301), .B(n30626), .Y(n33448) );
  AND2X2 U10012 ( .A(n23282), .B(n30626), .Y(n33429) );
  AND2X2 U10013 ( .A(n27252), .B(n32491), .Y(n32533) );
  AND2X2 U10014 ( .A(n29943), .B(n29330), .Y(n32480) );
  AND2X2 U10015 ( .A(n23285), .B(n32491), .Y(n33021) );
  INVX1 U10016 ( .A(n20806), .Y(n21435) );
  AND2X2 U10017 ( .A(n23290), .B(n32491), .Y(n32536) );
  AND2X2 U10018 ( .A(n23446), .B(n29331), .Y(n32477) );
  AND2X2 U10019 ( .A(n30626), .B(n23291), .Y(n33307) );
  AND2X2 U10020 ( .A(n23293), .B(n32491), .Y(n33002) );
  AND2X2 U10021 ( .A(n29993), .B(n29331), .Y(n32770) );
  AND2X2 U10022 ( .A(n30626), .B(n23294), .Y(n33276) );
  AND2X2 U10023 ( .A(n23295), .B(n32491), .Y(n32895) );
  AND2X2 U10024 ( .A(n30002), .B(n25723), .Y(n32478) );
  AND2X2 U10025 ( .A(n27268), .B(n25721), .Y(n31924) );
  AND2X2 U10026 ( .A(n21405), .B(n25720), .Y(n31929) );
  AND2X2 U10027 ( .A(n25721), .B(n23442), .Y(n31934) );
  AND2X2 U10028 ( .A(n27307), .B(n25721), .Y(n31939) );
  AND2X2 U10029 ( .A(n27308), .B(n25720), .Y(n31944) );
  AND2X2 U10030 ( .A(n27269), .B(n25720), .Y(n31949) );
  AND2X2 U10031 ( .A(n30410), .B(n25721), .Y(n31954) );
  AND2X2 U10032 ( .A(n27306), .B(n26163), .Y(n31960) );
  AND2X2 U10033 ( .A(n27306), .B(n27268), .Y(n31965) );
  AND2X2 U10034 ( .A(n27306), .B(n21405), .Y(n31970) );
  AND2X2 U10035 ( .A(n27306), .B(n27307), .Y(n31979) );
  AND2X2 U10036 ( .A(n27306), .B(n27308), .Y(n31984) );
  AND2X2 U10037 ( .A(n27306), .B(n27269), .Y(n31989) );
  AND2X2 U10038 ( .A(n27306), .B(n30410), .Y(n31995) );
  AND2X1 U10039 ( .A(n30226), .B(n27307), .Y(n32008) );
  AND2X2 U10040 ( .A(n30226), .B(n27269), .Y(n32014) );
  AND2X2 U10041 ( .A(n21414), .B(n26163), .Y(n32020) );
  AND2X2 U10042 ( .A(n21414), .B(n21405), .Y(n32026) );
  AND2X2 U10043 ( .A(n21414), .B(n27307), .Y(n32032) );
  AND2X2 U10044 ( .A(n21414), .B(n27269), .Y(n32038) );
  AND2X2 U10045 ( .A(n27266), .B(n26163), .Y(n32046) );
  AND2X2 U10046 ( .A(n27266), .B(n27268), .Y(n32050) );
  AND2X2 U10047 ( .A(n27266), .B(n21405), .Y(n32054) );
  AND2X2 U10048 ( .A(n27266), .B(n27307), .Y(n32061) );
  AND2X2 U10049 ( .A(n27266), .B(n27308), .Y(n32065) );
  AND2X2 U10050 ( .A(n27266), .B(n27269), .Y(n32069) );
  AND2X2 U10051 ( .A(n27266), .B(n30410), .Y(n32073) );
  AND2X2 U10052 ( .A(n27305), .B(n26163), .Y(n32077) );
  AND2X1 U10053 ( .A(n27305), .B(n27268), .Y(n32081) );
  AND2X2 U10054 ( .A(n27305), .B(n21405), .Y(n32085) );
  AND2X2 U10055 ( .A(n27305), .B(n27307), .Y(n32092) );
  AND2X2 U10056 ( .A(n27305), .B(n27308), .Y(n32096) );
  AND2X2 U10057 ( .A(n27305), .B(n27269), .Y(n32102) );
  AND2X2 U10058 ( .A(n27305), .B(n30410), .Y(n32106) );
  AND2X2 U10059 ( .A(n27264), .B(n26163), .Y(n32109) );
  AND2X2 U10060 ( .A(n30411), .B(n27237), .Y(n32112) );
  AND2X2 U10061 ( .A(n27264), .B(n21405), .Y(n32115) );
  AND2X2 U10062 ( .A(n27264), .B(n27307), .Y(n32121) );
  AND2X1 U10063 ( .A(n27264), .B(n27269), .Y(n32127) );
  AND2X2 U10064 ( .A(n29670), .B(n26163), .Y(n32132) );
  AND2X2 U10065 ( .A(n21405), .B(n29670), .Y(n32138) );
  AND2X2 U10066 ( .A(n27307), .B(n29670), .Y(n32144) );
  AND2X2 U10067 ( .A(n27269), .B(n29670), .Y(n32149) );
  AND2X2 U10068 ( .A(n30473), .B(n30472), .Y(n32154) );
  AND2X2 U10069 ( .A(n31868), .B(n22794), .Y(n31891) );
  AND2X1 U10070 ( .A(n30656), .B(net96340), .Y(n31876) );
  INVX1 U10071 ( .A(n31876), .Y(n21438) );
  AND2X2 U10072 ( .A(n25871), .B(n32234), .Y(n30823) );
  INVX1 U10073 ( .A(n30823), .Y(n21441) );
  AND2X2 U10074 ( .A(n25872), .B(n32239), .Y(n30844) );
  INVX1 U10075 ( .A(n30844), .Y(n21444) );
  AND2X2 U10076 ( .A(n27235), .B(n31868), .Y(n31897) );
  AND2X2 U10077 ( .A(n25886), .B(n32323), .Y(n31217) );
  INVX1 U10078 ( .A(n31217), .Y(n21447) );
  AND2X2 U10079 ( .A(n25882), .B(n32331), .Y(n31257) );
  INVX1 U10080 ( .A(n31257), .Y(n21450) );
  AND2X2 U10081 ( .A(n25880), .B(n32339), .Y(n31294) );
  INVX1 U10082 ( .A(n31294), .Y(n21453) );
  AND2X2 U10083 ( .A(n25876), .B(n32343), .Y(n31313) );
  INVX1 U10084 ( .A(n31313), .Y(n21456) );
  AND2X2 U10085 ( .A(n25879), .B(n32347), .Y(n31331) );
  INVX1 U10086 ( .A(n31331), .Y(n21459) );
  AND2X2 U10087 ( .A(n25884), .B(n32351), .Y(n31351) );
  INVX1 U10088 ( .A(n31351), .Y(n21462) );
  AND2X2 U10089 ( .A(n25870), .B(n32355), .Y(n31371) );
  INVX1 U10090 ( .A(n31371), .Y(n21465) );
  AND2X2 U10091 ( .A(n25881), .B(n32359), .Y(n31391) );
  INVX1 U10092 ( .A(n31391), .Y(n21467) );
  AND2X2 U10093 ( .A(n25878), .B(n32363), .Y(n31411) );
  INVX1 U10094 ( .A(n31411), .Y(n21469) );
  AND2X2 U10095 ( .A(n25877), .B(n32367), .Y(n31432) );
  INVX1 U10096 ( .A(n31432), .Y(n21472) );
  AND2X2 U10097 ( .A(n25930), .B(n32371), .Y(n31451) );
  INVX1 U10098 ( .A(n31451), .Y(n21475) );
  AND2X2 U10099 ( .A(n25929), .B(n32375), .Y(n31471) );
  INVX1 U10100 ( .A(n31471), .Y(n21478) );
  AND2X2 U10101 ( .A(n25916), .B(n32379), .Y(n31490) );
  INVX1 U10102 ( .A(n31490), .Y(n21481) );
  AND2X2 U10103 ( .A(n25931), .B(n32383), .Y(n31509) );
  INVX1 U10104 ( .A(n31509), .Y(n21484) );
  AND2X2 U10105 ( .A(n29378), .B(n31600), .Y(n31612) );
  INVX1 U10106 ( .A(n31612), .Y(n21487) );
  AND2X2 U10107 ( .A(n29376), .B(n31637), .Y(n31648) );
  AND2X2 U10108 ( .A(net109585), .B(net96340), .Y(n34174) );
  AND2X2 U10109 ( .A(n3260), .B(n23451), .Y(n32482) );
  INVX1 U10110 ( .A(n32482), .Y(n21490) );
  AND2X2 U10111 ( .A(n3194), .B(n23471), .Y(n32493) );
  INVX1 U10112 ( .A(n32493), .Y(n21493) );
  AND2X2 U10113 ( .A(n3152), .B(n21212), .Y(n32503) );
  AND2X2 U10114 ( .A(n3208), .B(n32528), .Y(n32531) );
  INVX1 U10115 ( .A(n32531), .Y(n21496) );
  AND2X2 U10116 ( .A(n3180), .B(n32783), .Y(n32590) );
  AND2X2 U10117 ( .A(n3150), .B(n32792), .Y(n32599) );
  AND2X2 U10118 ( .A(n3178), .B(n33609), .Y(n32643) );
  INVX1 U10119 ( .A(n32643), .Y(n21499) );
  AND2X2 U10120 ( .A(n3274), .B(n32764), .Y(n32672) );
  INVX1 U10121 ( .A(n32672), .Y(n21502) );
  AND2X2 U10122 ( .A(n32777), .B(n3208), .Y(n32682) );
  AND2X2 U10123 ( .A(n3160), .B(n27232), .Y(n32691) );
  AND2X2 U10124 ( .A(n3210), .B(n32528), .Y(n32719) );
  INVX1 U10125 ( .A(n32719), .Y(n21505) );
  AND2X2 U10126 ( .A(n3248), .B(n33326), .Y(n32729) );
  AND2X2 U10127 ( .A(n3182), .B(n33609), .Y(n32737) );
  AND2X2 U10128 ( .A(n29331), .B(n21221), .Y(n32779) );
  AND2X2 U10129 ( .A(n3161), .B(n27232), .Y(n32788) );
  AND2X2 U10130 ( .A(n33326), .B(n3249), .Y(n32825) );
  INVX1 U10131 ( .A(n32825), .Y(n21508) );
  AND2X2 U10132 ( .A(n33609), .B(n3183), .Y(n32833) );
  AND2X2 U10133 ( .A(n3195), .B(n32489), .Y(n32868) );
  AND2X2 U10134 ( .A(n32792), .B(n3153), .Y(n32879) );
  INVX1 U10135 ( .A(n32918), .Y(n21511) );
  AND2X2 U10136 ( .A(n3245), .B(n33326), .Y(n33026) );
  AND2X2 U10137 ( .A(n3179), .B(n33609), .Y(n33035) );
  INVX1 U10138 ( .A(n33035), .Y(n21514) );
  AND2X2 U10139 ( .A(n23068), .B(n22089), .Y(n33073) );
  OR2X2 U10140 ( .A(n33095), .B(n33103), .Y(n33102) );
  INVX1 U10141 ( .A(n33102), .Y(n21517) );
  AND2X2 U10142 ( .A(T[1]), .B(n25111), .Y(n33122) );
  AND2X2 U10143 ( .A(T[3]), .B(n25650), .Y(n33128) );
  AND2X2 U10144 ( .A(n34360), .B(n25621), .Y(n33132) );
  AND2X2 U10145 ( .A(n25339), .B(n25419), .Y(n33157) );
  OR2X2 U10146 ( .A(n33131), .B(n33130), .Y(n33139) );
  INVX1 U10147 ( .A(n33139), .Y(n21520) );
  AND2X2 U10148 ( .A(n25337), .B(n33133), .Y(n33135) );
  INVX1 U10149 ( .A(n33135), .Y(n21522) );
  AND2X2 U10150 ( .A(T[4]), .B(n34232), .Y(n34246) );
  AND2X2 U10151 ( .A(n34356), .B(n34233), .Y(n34243) );
  AND2X2 U10152 ( .A(n34323), .B(n34249), .Y(n34257) );
  INVX1 U10153 ( .A(n34257), .Y(n21523) );
  AND2X2 U10154 ( .A(n25761), .B(n34309), .Y(n34261) );
  AND2X2 U10155 ( .A(n34317), .B(n25159), .Y(n34259) );
  AND2X2 U10156 ( .A(n34417), .B(n34263), .Y(n34272) );
  INVX1 U10157 ( .A(n34272), .Y(n21524) );
  AND2X2 U10158 ( .A(T[3]), .B(n23919), .Y(n34303) );
  AND2X2 U10159 ( .A(n23072), .B(n25446), .Y(n34324) );
  AND2X2 U10160 ( .A(n25664), .B(n25405), .Y(n34401) );
  INVX1 U10161 ( .A(n34401), .Y(n21525) );
  BUFX2 U10162 ( .A(n29483), .Y(n21526) );
  BUFX2 U10163 ( .A(n29578), .Y(n21527) );
  BUFX2 U10164 ( .A(n32541), .Y(n21528) );
  BUFX2 U10165 ( .A(n32632), .Y(n21529) );
  BUFX2 U10166 ( .A(n32824), .Y(n21530) );
  BUFX2 U10167 ( .A(n32926), .Y(n21531) );
  BUFX2 U10168 ( .A(n33034), .Y(n21532) );
  BUFX2 U10169 ( .A(n33975), .Y(n21533) );
  BUFX2 U10170 ( .A(n33977), .Y(n21534) );
  BUFX2 U10171 ( .A(n33981), .Y(n21535) );
  BUFX2 U10172 ( .A(n33987), .Y(n21536) );
  BUFX2 U10173 ( .A(n34181), .Y(n21537) );
  BUFX2 U10174 ( .A(n34201), .Y(n21538) );
  BUFX2 U10175 ( .A(n34217), .Y(n21539) );
  BUFX2 U10176 ( .A(n34289), .Y(n21540) );
  BUFX2 U10177 ( .A(n34348), .Y(n21541) );
  AND2X2 U10178 ( .A(n25475), .B(n29197), .Y(n25476) );
  INVX1 U10179 ( .A(n25476), .Y(n21542) );
  AND2X2 U10180 ( .A(n27281), .B(n33386), .Y(n25520) );
  INVX1 U10181 ( .A(n25520), .Y(n21543) );
  AND2X2 U10182 ( .A(n27220), .B(n3129), .Y(n25586) );
  INVX1 U10183 ( .A(n25586), .Y(n21544) );
  AND2X2 U10184 ( .A(n3167), .B(n26519), .Y(n27141) );
  INVX1 U10185 ( .A(n27141), .Y(n21545) );
  AND2X2 U10186 ( .A(n33726), .B(n3145), .Y(n27144) );
  INVX1 U10187 ( .A(n27144), .Y(n21546) );
  BUFX2 U10188 ( .A(n32802), .Y(n21547) );
  BUFX2 U10189 ( .A(n33201), .Y(n21548) );
  BUFX2 U10190 ( .A(n33231), .Y(n21549) );
  BUFX2 U10191 ( .A(n33384), .Y(n21550) );
  BUFX2 U10192 ( .A(n34186), .Y(n21551) );
  BUFX2 U10193 ( .A(n34205), .Y(n21552) );
  AND2X2 U10194 ( .A(n24004), .B(n22025), .Y(n30935) );
  INVX1 U10195 ( .A(n30935), .Y(n21553) );
  AND2X2 U10196 ( .A(n25519), .B(n22039), .Y(n31152) );
  INVX1 U10197 ( .A(n31152), .Y(n21554) );
  AND2X2 U10198 ( .A(n27216), .B(n3117), .Y(n25587) );
  INVX1 U10199 ( .A(n25587), .Y(n21555) );
  INVX1 U10200 ( .A(n25343), .Y(n21556) );
  AND2X2 U10201 ( .A(direction_lee[2]), .B(n21210), .Y(n29488) );
  INVX1 U10202 ( .A(n29488), .Y(n21557) );
  AND2X2 U10203 ( .A(n23947), .B(n21080), .Y(n31896) );
  INVX1 U10204 ( .A(n31896), .Y(n21558) );
  INVX1 U10205 ( .A(n25706), .Y(n21559) );
  INVX1 U10206 ( .A(n25726), .Y(n21560) );
  BUFX2 U10207 ( .A(n29474), .Y(n21561) );
  BUFX2 U10208 ( .A(n29495), .Y(n21562) );
  BUFX2 U10209 ( .A(n29497), .Y(n21563) );
  BUFX2 U10210 ( .A(n29568), .Y(n21564) );
  BUFX2 U10211 ( .A(n29574), .Y(n21565) );
  BUFX2 U10212 ( .A(n29576), .Y(n21566) );
  BUFX2 U10213 ( .A(n32158), .Y(n21567) );
  BUFX2 U10214 ( .A(n32163), .Y(n21568) );
  BUFX2 U10215 ( .A(n32168), .Y(n21569) );
  BUFX2 U10216 ( .A(n32173), .Y(n21570) );
  BUFX2 U10217 ( .A(n32178), .Y(n21571) );
  BUFX2 U10218 ( .A(n32183), .Y(n21572) );
  BUFX2 U10219 ( .A(n32466), .Y(n21573) );
  BUFX2 U10220 ( .A(n32467), .Y(n21574) );
  BUFX2 U10221 ( .A(n32471), .Y(n21575) );
  BUFX2 U10222 ( .A(n32473), .Y(n21576) );
  BUFX2 U10223 ( .A(n32484), .Y(n21577) );
  BUFX2 U10224 ( .A(n32485), .Y(n21578) );
  BUFX2 U10225 ( .A(n32495), .Y(n21579) );
  BUFX2 U10226 ( .A(n32497), .Y(n21580) );
  BUFX2 U10227 ( .A(n32505), .Y(n21581) );
  BUFX2 U10228 ( .A(n32507), .Y(n21582) );
  BUFX2 U10229 ( .A(n32516), .Y(n21583) );
  BUFX2 U10230 ( .A(n32519), .Y(n21584) );
  BUFX2 U10231 ( .A(n32522), .Y(n21585) );
  BUFX2 U10232 ( .A(n32524), .Y(n21586) );
  BUFX2 U10233 ( .A(n32534), .Y(n21587) );
  BUFX2 U10234 ( .A(n32537), .Y(n21588) );
  BUFX2 U10235 ( .A(n32544), .Y(n21589) );
  BUFX2 U10236 ( .A(n32545), .Y(n21590) );
  BUFX2 U10237 ( .A(n32554), .Y(n21591) );
  BUFX2 U10238 ( .A(n32555), .Y(n21592) );
  BUFX2 U10239 ( .A(n32566), .Y(n21593) );
  BUFX2 U10240 ( .A(n32568), .Y(n21594) );
  BUFX2 U10241 ( .A(n32572), .Y(n21595) );
  BUFX2 U10242 ( .A(n32574), .Y(n21596) );
  BUFX2 U10243 ( .A(n32581), .Y(n21597) );
  BUFX2 U10244 ( .A(n32583), .Y(n21598) );
  BUFX2 U10245 ( .A(n32592), .Y(n21666) );
  BUFX2 U10246 ( .A(n32594), .Y(n21699) );
  BUFX2 U10247 ( .A(n32601), .Y(n21767) );
  BUFX2 U10248 ( .A(n32603), .Y(n21782) );
  BUFX2 U10249 ( .A(n32613), .Y(n21801) );
  BUFX2 U10250 ( .A(n32614), .Y(n21848) );
  BUFX2 U10251 ( .A(n32617), .Y(n21849) );
  BUFX2 U10252 ( .A(n32618), .Y(n21850) );
  BUFX2 U10253 ( .A(n32626), .Y(n21851) );
  BUFX2 U10254 ( .A(n32637), .Y(n21853) );
  BUFX2 U10255 ( .A(n32645), .Y(n21855) );
  BUFX2 U10256 ( .A(n32647), .Y(n21856) );
  BUFX2 U10257 ( .A(n32658), .Y(n21857) );
  BUFX2 U10258 ( .A(n32660), .Y(n21859) );
  BUFX2 U10259 ( .A(n32664), .Y(n21861) );
  BUFX2 U10260 ( .A(n32666), .Y(n21862) );
  BUFX2 U10261 ( .A(n32674), .Y(n21863) );
  BUFX2 U10262 ( .A(n32676), .Y(n21864) );
  BUFX2 U10263 ( .A(n32684), .Y(n21865) );
  BUFX2 U10264 ( .A(n32686), .Y(n21866) );
  BUFX2 U10265 ( .A(n32693), .Y(n21867) );
  BUFX2 U10266 ( .A(n32695), .Y(n21868) );
  BUFX2 U10267 ( .A(n32705), .Y(n21869) );
  BUFX2 U10268 ( .A(n32707), .Y(n21870) );
  BUFX2 U10269 ( .A(n32711), .Y(n21871) );
  BUFX2 U10270 ( .A(n32721), .Y(n21872) );
  BUFX2 U10271 ( .A(n32731), .Y(n21873) );
  BUFX2 U10272 ( .A(n32732), .Y(n21874) );
  BUFX2 U10273 ( .A(n32739), .Y(n21875) );
  BUFX2 U10274 ( .A(n32741), .Y(n21876) );
  BUFX2 U10275 ( .A(n32752), .Y(n21877) );
  BUFX2 U10276 ( .A(n32753), .Y(n21878) );
  BUFX2 U10277 ( .A(n32757), .Y(n21879) );
  BUFX2 U10278 ( .A(n32759), .Y(n21880) );
  BUFX2 U10279 ( .A(n32768), .Y(n21881) );
  BUFX2 U10280 ( .A(n32771), .Y(n21882) );
  BUFX2 U10281 ( .A(n32781), .Y(n21883) );
  BUFX2 U10282 ( .A(n32784), .Y(n21884) );
  BUFX2 U10283 ( .A(n32790), .Y(n21885) );
  BUFX2 U10284 ( .A(n32793), .Y(n21886) );
  BUFX2 U10285 ( .A(n32804), .Y(n21887) );
  BUFX2 U10286 ( .A(n32808), .Y(n21888) );
  BUFX2 U10287 ( .A(n32810), .Y(n21889) );
  BUFX2 U10288 ( .A(n32818), .Y(n21890) );
  BUFX2 U10289 ( .A(n32819), .Y(n21891) );
  BUFX2 U10290 ( .A(n32827), .Y(n21892) );
  BUFX2 U10291 ( .A(n32828), .Y(n21893) );
  BUFX2 U10292 ( .A(n32835), .Y(n21894) );
  BUFX2 U10293 ( .A(n32836), .Y(n21895) );
  BUFX2 U10294 ( .A(n32847), .Y(n21896) );
  BUFX2 U10295 ( .A(n32849), .Y(n21897) );
  BUFX2 U10296 ( .A(n32862), .Y(n21898) );
  BUFX2 U10297 ( .A(n32864), .Y(n21899) );
  BUFX2 U10298 ( .A(n32870), .Y(n21900) );
  BUFX2 U10299 ( .A(n32873), .Y(n21901) );
  BUFX2 U10300 ( .A(n32881), .Y(n21902) );
  BUFX2 U10301 ( .A(n32893), .Y(n21903) );
  BUFX2 U10302 ( .A(n32896), .Y(n21904) );
  BUFX2 U10303 ( .A(n32900), .Y(n21905) );
  BUFX2 U10304 ( .A(n32911), .Y(n21906) );
  BUFX2 U10305 ( .A(n32920), .Y(n21907) );
  BUFX2 U10306 ( .A(n32921), .Y(n21908) );
  BUFX2 U10307 ( .A(n32929), .Y(n21909) );
  BUFX2 U10308 ( .A(n32941), .Y(n21910) );
  BUFX2 U10309 ( .A(n32943), .Y(n21911) );
  BUFX2 U10310 ( .A(n32948), .Y(n21912) );
  BUFX2 U10311 ( .A(n32962), .Y(n21913) );
  BUFX2 U10312 ( .A(n32965), .Y(n21914) );
  BUFX2 U10313 ( .A(n32976), .Y(n21915) );
  BUFX2 U10314 ( .A(n32979), .Y(n21916) );
  BUFX2 U10315 ( .A(n32986), .Y(n21917) );
  BUFX2 U10316 ( .A(n32989), .Y(n21918) );
  BUFX2 U10317 ( .A(n33001), .Y(n21919) );
  BUFX2 U10318 ( .A(n33003), .Y(n21920) );
  BUFX2 U10319 ( .A(n33009), .Y(n21921) );
  BUFX2 U10320 ( .A(n33028), .Y(n21922) );
  BUFX2 U10321 ( .A(n33030), .Y(n21923) );
  BUFX2 U10322 ( .A(n34212), .Y(n21924) );
  BUFX2 U10323 ( .A(n34274), .Y(n21925) );
  BUFX2 U10324 ( .A(n30640), .Y(n21926) );
  BUFX2 U10325 ( .A(n30671), .Y(n21927) );
  BUFX2 U10326 ( .A(n30694), .Y(n21928) );
  BUFX2 U10327 ( .A(n30714), .Y(n21929) );
  BUFX2 U10328 ( .A(n30733), .Y(n21930) );
  BUFX2 U10329 ( .A(n30773), .Y(n21931) );
  BUFX2 U10330 ( .A(n30794), .Y(n21932) );
  BUFX2 U10331 ( .A(n30813), .Y(n21933) );
  BUFX2 U10332 ( .A(n30834), .Y(n21934) );
  BUFX2 U10333 ( .A(n30853), .Y(n21935) );
  BUFX2 U10334 ( .A(n30915), .Y(n21936) );
  BUFX2 U10335 ( .A(n30955), .Y(n21937) );
  BUFX2 U10336 ( .A(n30976), .Y(n21938) );
  BUFX2 U10337 ( .A(n31012), .Y(n21939) );
  BUFX2 U10338 ( .A(n31033), .Y(n21940) );
  BUFX2 U10339 ( .A(n31071), .Y(n21941) );
  BUFX2 U10340 ( .A(n31090), .Y(n21942) );
  BUFX2 U10341 ( .A(n31111), .Y(n21943) );
  BUFX2 U10342 ( .A(n31130), .Y(n21944) );
  BUFX2 U10343 ( .A(n31188), .Y(n21945) );
  BUFX2 U10344 ( .A(n31207), .Y(n21946) );
  BUFX2 U10345 ( .A(n31228), .Y(n21947) );
  BUFX2 U10346 ( .A(n31247), .Y(n21948) );
  BUFX2 U10347 ( .A(n31268), .Y(n21949) );
  BUFX2 U10348 ( .A(n31285), .Y(n21950) );
  BUFX2 U10349 ( .A(n31321), .Y(n21951) );
  BUFX2 U10350 ( .A(n31361), .Y(n21952) );
  BUFX2 U10351 ( .A(n31381), .Y(n21953) );
  BUFX2 U10352 ( .A(n31401), .Y(n21954) );
  BUFX2 U10353 ( .A(n31461), .Y(n21955) );
  BUFX2 U10354 ( .A(n31481), .Y(n21956) );
  BUFX2 U10355 ( .A(n31518), .Y(n21957) );
  BUFX2 U10356 ( .A(n31538), .Y(n21958) );
  BUFX2 U10357 ( .A(n31558), .Y(n21959) );
  BUFX2 U10358 ( .A(n31599), .Y(n21960) );
  BUFX2 U10359 ( .A(n31619), .Y(n21961) );
  BUFX2 U10360 ( .A(n31655), .Y(n21962) );
  BUFX2 U10361 ( .A(n31673), .Y(n21963) );
  BUFX2 U10362 ( .A(n31693), .Y(n21964) );
  BUFX2 U10363 ( .A(n31712), .Y(n21965) );
  BUFX2 U10364 ( .A(n31733), .Y(n21966) );
  BUFX2 U10365 ( .A(n31750), .Y(n21967) );
  BUFX2 U10366 ( .A(n31771), .Y(n21968) );
  BUFX2 U10367 ( .A(n31810), .Y(n21969) );
  BUFX2 U10368 ( .A(n31829), .Y(n21970) );
  BUFX2 U10369 ( .A(n33184), .Y(n21971) );
  BUFX2 U10370 ( .A(n33210), .Y(n21972) );
  BUFX2 U10371 ( .A(n33219), .Y(n21973) );
  BUFX2 U10372 ( .A(n33241), .Y(n21974) );
  BUFX2 U10373 ( .A(n33250), .Y(n21975) );
  BUFX2 U10374 ( .A(n33271), .Y(n21976) );
  BUFX2 U10375 ( .A(n33280), .Y(n21977) );
  BUFX2 U10376 ( .A(n33302), .Y(n21978) );
  BUFX2 U10377 ( .A(n33311), .Y(n21979) );
  BUFX2 U10378 ( .A(n33333), .Y(n21980) );
  BUFX2 U10379 ( .A(n33342), .Y(n21981) );
  BUFX2 U10380 ( .A(n33363), .Y(n21982) );
  BUFX2 U10381 ( .A(n33393), .Y(n21983) );
  BUFX2 U10382 ( .A(n33402), .Y(n21984) );
  BUFX2 U10383 ( .A(n33424), .Y(n21985) );
  BUFX2 U10384 ( .A(n34258), .Y(n21986) );
  BUFX2 U10385 ( .A(n34377), .Y(n21987) );
  INVX1 U10386 ( .A(n25213), .Y(n21988) );
  OR2X2 U10387 ( .A(n25474), .B(n29194), .Y(n30874) );
  INVX1 U10388 ( .A(n30874), .Y(n21989) );
  OR2X2 U10389 ( .A(n21357), .B(n26285), .Y(n31168) );
  INVX1 U10390 ( .A(n31168), .Y(n21990) );
  AND2X2 U10391 ( .A(n32191), .B(n27263), .Y(n32192) );
  INVX1 U10392 ( .A(n32192), .Y(n21991) );
  INVX1 U10393 ( .A(n25697), .Y(n21992) );
  INVX1 U10394 ( .A(n34269), .Y(n21993) );
  BUFX2 U10395 ( .A(n29588), .Y(n21994) );
  BUFX2 U10396 ( .A(n32161), .Y(n21995) );
  BUFX2 U10397 ( .A(n33434), .Y(n21996) );
  BUFX2 U10398 ( .A(n33681), .Y(n21997) );
  BUFX2 U10399 ( .A(n33686), .Y(n21998) );
  BUFX2 U10400 ( .A(n33703), .Y(n21999) );
  BUFX2 U10401 ( .A(n33725), .Y(n22000) );
  BUFX2 U10402 ( .A(n33730), .Y(n22001) );
  BUFX2 U10403 ( .A(n33746), .Y(n22002) );
  BUFX2 U10404 ( .A(n33752), .Y(n22003) );
  BUFX2 U10405 ( .A(n33769), .Y(n22004) );
  BUFX2 U10406 ( .A(n33774), .Y(n22005) );
  BUFX2 U10407 ( .A(n33791), .Y(n22006) );
  BUFX2 U10408 ( .A(n33796), .Y(n22007) );
  BUFX2 U10409 ( .A(n33813), .Y(n22008) );
  BUFX2 U10410 ( .A(n33819), .Y(n22009) );
  BUFX2 U10411 ( .A(n33836), .Y(n22010) );
  BUFX2 U10412 ( .A(n33841), .Y(n22011) );
  BUFX2 U10413 ( .A(n33859), .Y(n22012) );
  BUFX2 U10414 ( .A(n33865), .Y(n22013) );
  BUFX2 U10415 ( .A(n33882), .Y(n22014) );
  BUFX2 U10416 ( .A(n33889), .Y(n22015) );
  BUFX2 U10417 ( .A(n33925), .Y(n22016) );
  BUFX2 U10418 ( .A(n33940), .Y(n22017) );
  BUFX2 U10419 ( .A(n33948), .Y(n22018) );
  BUFX2 U10420 ( .A(n33950), .Y(n22019) );
  BUFX2 U10421 ( .A(n33956), .Y(n22020) );
  BUFX2 U10422 ( .A(n33966), .Y(n22021) );
  BUFX2 U10423 ( .A(n33985), .Y(n22022) );
  BUFX2 U10424 ( .A(n33991), .Y(n22023) );
  BUFX2 U10425 ( .A(n34191), .Y(n22024) );
  BUFX2 U10426 ( .A(n30934), .Y(n22025) );
  BUFX2 U10427 ( .A(n33447), .Y(n22026) );
  BUFX2 U10428 ( .A(n33492), .Y(n22027) );
  BUFX2 U10429 ( .A(n33498), .Y(n22028) );
  BUFX2 U10430 ( .A(n33515), .Y(n22029) );
  BUFX2 U10431 ( .A(n33571), .Y(n22030) );
  BUFX2 U10432 ( .A(n33577), .Y(n22031) );
  BUFX2 U10433 ( .A(n33594), .Y(n22032) );
  BUFX2 U10434 ( .A(n33599), .Y(n22033) );
  BUFX2 U10435 ( .A(n33621), .Y(n22034) );
  BUFX2 U10436 ( .A(n33637), .Y(n22035) );
  BUFX2 U10437 ( .A(n33643), .Y(n22036) );
  BUFX2 U10438 ( .A(n33660), .Y(n22037) );
  BUFX2 U10439 ( .A(n33665), .Y(n22038) );
  OR2X2 U10440 ( .A(n25518), .B(n26279), .Y(n31151) );
  INVX1 U10441 ( .A(n31151), .Y(n22039) );
  AND2X2 U10442 ( .A(direction_lee[0]), .B(n21125), .Y(n29487) );
  AND2X2 U10443 ( .A(n33609), .B(n3181), .Y(n32927) );
  INVX1 U10444 ( .A(n32927), .Y(n22040) );
  BUFX2 U10445 ( .A(n29589), .Y(n22041) );
  BUFX2 U10446 ( .A(n32826), .Y(n22042) );
  BUFX2 U10447 ( .A(n32928), .Y(n22043) );
  BUFX2 U10448 ( .A(n33036), .Y(n22044) );
  BUFX2 U10449 ( .A(n33936), .Y(n22045) );
  BUFX2 U10450 ( .A(n33938), .Y(n22046) );
  BUFX2 U10451 ( .A(n33942), .Y(n22047) );
  BUFX2 U10452 ( .A(n33944), .Y(n22048) );
  BUFX2 U10453 ( .A(n33946), .Y(n22049) );
  BUFX2 U10454 ( .A(n33952), .Y(n22050) );
  BUFX2 U10455 ( .A(n33954), .Y(n22051) );
  BUFX2 U10456 ( .A(n33958), .Y(n22052) );
  BUFX2 U10457 ( .A(n33960), .Y(n22057) );
  BUFX2 U10458 ( .A(n33962), .Y(n22061) );
  BUFX2 U10459 ( .A(n33964), .Y(n22062) );
  BUFX2 U10460 ( .A(n33968), .Y(n22065) );
  BUFX2 U10461 ( .A(n33970), .Y(n22069) );
  BUFX2 U10462 ( .A(net90010), .Y(net144199) );
  BUFX2 U10463 ( .A(n33973), .Y(n22070) );
  BUFX2 U10464 ( .A(n33979), .Y(n22073) );
  BUFX2 U10465 ( .A(n33983), .Y(n22077) );
  BUFX2 U10466 ( .A(n33989), .Y(n22078) );
  BUFX2 U10467 ( .A(n34184), .Y(n22081) );
  BUFX2 U10468 ( .A(n34268), .Y(n22085) );
  AND2X2 U10469 ( .A(n3185), .B(n33019), .Y(n27043) );
  INVX1 U10470 ( .A(n27043), .Y(n22086) );
  INVX1 U10471 ( .A(n25767), .Y(n22089) );
  BUFX2 U10472 ( .A(n34339), .Y(n22094) );
  AND2X2 U10473 ( .A(n21542), .B(n26971), .Y(n31779) );
  INVX1 U10474 ( .A(n31779), .Y(n22097) );
  BUFX2 U10475 ( .A(n31915), .Y(n22102) );
  BUFX2 U10476 ( .A(n29535), .Y(n22109) );
  BUFX2 U10477 ( .A(n29721), .Y(n22110) );
  BUFX2 U10478 ( .A(n29717), .Y(n22113) );
  AND2X2 U10479 ( .A(n25572), .B(n21547), .Y(n32807) );
  INVX1 U10480 ( .A(n32807), .Y(n22118) );
  BUFX2 U10481 ( .A(n33181), .Y(n22122) );
  BUFX2 U10482 ( .A(n33191), .Y(n22126) );
  BUFX2 U10483 ( .A(n29534), .Y(n22129) );
  BUFX2 U10484 ( .A(n29709), .Y(n22130) );
  BUFX2 U10485 ( .A(n29716), .Y(n22134) );
  INVX1 U10486 ( .A(n29720), .Y(n22138) );
  AND2X2 U10487 ( .A(n29550), .B(n26697), .Y(n29551) );
  INVX1 U10488 ( .A(n29551), .Y(n22142) );
  BUFX2 U10489 ( .A(n29554), .Y(n22145) );
  BUFX2 U10490 ( .A(n34416), .Y(n22146) );
  AND2X2 U10491 ( .A(n23076), .B(n25224), .Y(n30646) );
  INVX1 U10492 ( .A(n30646), .Y(n22150) );
  AND2X2 U10493 ( .A(n23189), .B(n23146), .Y(n30674) );
  INVX1 U10494 ( .A(n30674), .Y(n22154) );
  AND2X2 U10495 ( .A(n25184), .B(n23148), .Y(n30697) );
  INVX1 U10496 ( .A(n30697), .Y(n22158) );
  AND2X2 U10497 ( .A(n25185), .B(n23149), .Y(n30717) );
  INVX1 U10498 ( .A(n30717), .Y(n22162) );
  AND2X2 U10499 ( .A(n25186), .B(n23150), .Y(n30736) );
  INVX1 U10500 ( .A(n30736), .Y(n22166) );
  AND2X2 U10501 ( .A(n25187), .B(n23152), .Y(n30757) );
  INVX1 U10502 ( .A(n30757), .Y(n22169) );
  AND2X2 U10503 ( .A(n25188), .B(n23154), .Y(n30776) );
  INVX1 U10504 ( .A(n30776), .Y(n22170) );
  AND2X2 U10505 ( .A(n25189), .B(n23156), .Y(n30816) );
  INVX1 U10506 ( .A(n30816), .Y(n22174) );
  AND2X2 U10507 ( .A(n23190), .B(n23008), .Y(n30837) );
  INVX1 U10508 ( .A(n30837), .Y(n22177) );
  AND2X2 U10509 ( .A(n23192), .B(n23157), .Y(n30856) );
  INVX1 U10510 ( .A(n30856), .Y(n22178) );
  AND2X2 U10511 ( .A(n23078), .B(n23009), .Y(n30877) );
  INVX1 U10512 ( .A(n30877), .Y(n22182) );
  AND2X2 U10513 ( .A(n23194), .B(n25172), .Y(n30937) );
  INVX1 U10514 ( .A(n30937), .Y(n22190) );
  AND2X2 U10515 ( .A(n23079), .B(n23014), .Y(n30979) );
  INVX1 U10516 ( .A(n30979), .Y(n22198) );
  AND2X2 U10517 ( .A(n23195), .B(n23159), .Y(n31015) );
  INVX1 U10518 ( .A(n31015), .Y(n22206) );
  AND2X2 U10519 ( .A(n23161), .B(n25190), .Y(n31053) );
  INVX1 U10520 ( .A(n31053), .Y(n22214) );
  AND2X2 U10521 ( .A(n23196), .B(n23163), .Y(n31093) );
  INVX1 U10522 ( .A(n31093), .Y(n22222) );
  AND2X2 U10523 ( .A(n23090), .B(n25175), .Y(n31171) );
  INVX1 U10524 ( .A(n31171), .Y(n22229) );
  AND2X2 U10525 ( .A(n25176), .B(n23165), .Y(n31210) );
  INVX1 U10526 ( .A(n31210), .Y(n22230) );
  AND2X2 U10527 ( .A(n25177), .B(n23167), .Y(n31250) );
  INVX1 U10528 ( .A(n31250), .Y(n22237) );
  AND2X2 U10529 ( .A(n23197), .B(n23036), .Y(n31324) );
  INVX1 U10530 ( .A(n31324), .Y(n22238) );
  AND2X2 U10531 ( .A(n25191), .B(n23169), .Y(n31404) );
  INVX1 U10532 ( .A(n31404), .Y(n22241) );
  AND2X2 U10533 ( .A(n23171), .B(n25192), .Y(n31425) );
  INVX1 U10534 ( .A(n31425), .Y(n22245) );
  AND2X2 U10535 ( .A(n23173), .B(n23042), .Y(n31445) );
  INVX1 U10536 ( .A(n31445), .Y(n22246) );
  AND2X2 U10537 ( .A(n23175), .B(n23044), .Y(n31521) );
  INVX1 U10538 ( .A(n31521), .Y(n22250) );
  AND2X2 U10539 ( .A(n23472), .B(n23177), .Y(n31541) );
  INVX1 U10540 ( .A(n31541), .Y(n22254) );
  AND2X2 U10541 ( .A(n23199), .B(n23179), .Y(n31561) );
  INVX1 U10542 ( .A(n31561), .Y(n22258) );
  AND2X2 U10543 ( .A(n23053), .B(n23180), .Y(n31676) );
  INVX1 U10544 ( .A(n31676), .Y(n22262) );
  AND2X2 U10545 ( .A(n23182), .B(n22999), .Y(n31715) );
  INVX1 U10546 ( .A(n31715), .Y(n22265) );
  AND2X2 U10547 ( .A(n25193), .B(n23184), .Y(n31753) );
  INVX1 U10548 ( .A(n31753), .Y(n22266) );
  AND2X2 U10549 ( .A(n23210), .B(n23186), .Y(n31872) );
  INVX1 U10550 ( .A(n31872), .Y(n22270) );
  AND2X2 U10551 ( .A(n33097), .B(n25167), .Y(n33098) );
  INVX1 U10552 ( .A(n33098), .Y(n22273) );
  AND2X2 U10553 ( .A(n33169), .B(n33168), .Y(n33170) );
  AND2X2 U10554 ( .A(n20952), .B(n25183), .Y(n34245) );
  INVX1 U10555 ( .A(n34245), .Y(n22274) );
  AND2X2 U10556 ( .A(n25642), .B(n25629), .Y(n34296) );
  INVX1 U10557 ( .A(n34296), .Y(n22278) );
  BUFX2 U10558 ( .A(n29597), .Y(n22282) );
  BUFX2 U10559 ( .A(n30682), .Y(n22286) );
  BUFX2 U10560 ( .A(n30845), .Y(n22290) );
  BUFX2 U10561 ( .A(n30864), .Y(n22294) );
  BUFX2 U10562 ( .A(n30880), .Y(n22298) );
  BUFX2 U10563 ( .A(n30885), .Y(n22302) );
  BUFX2 U10564 ( .A(n30905), .Y(n22306) );
  BUFX2 U10565 ( .A(n30926), .Y(n22307) );
  BUFX2 U10566 ( .A(n30945), .Y(n22310) );
  BUFX2 U10567 ( .A(n30966), .Y(n22311) );
  BUFX2 U10568 ( .A(n30982), .Y(n22312) );
  BUFX2 U10569 ( .A(n30986), .Y(n22313) );
  BUFX2 U10570 ( .A(n31000), .Y(n22314) );
  BUFX2 U10571 ( .A(n31023), .Y(n22315) );
  BUFX2 U10572 ( .A(n31037), .Y(n22316) );
  BUFX2 U10573 ( .A(n31061), .Y(n22317) );
  BUFX2 U10574 ( .A(n31075), .Y(n22318) );
  BUFX2 U10575 ( .A(n31082), .Y(n22319) );
  BUFX2 U10576 ( .A(n31101), .Y(n22320) );
  BUFX2 U10577 ( .A(n31115), .Y(n22321) );
  BUFX2 U10578 ( .A(n31122), .Y(n22322) );
  BUFX2 U10579 ( .A(n31141), .Y(n22375) );
  BUFX2 U10580 ( .A(n31155), .Y(n22420) );
  BUFX2 U10581 ( .A(n31178), .Y(n22421) );
  BUFX2 U10582 ( .A(n31192), .Y(n22422) );
  BUFX2 U10583 ( .A(n31199), .Y(n22423) );
  BUFX2 U10584 ( .A(n31232), .Y(n22424) );
  BUFX2 U10585 ( .A(n31272), .Y(n22434) );
  BUFX2 U10586 ( .A(n31295), .Y(n22437) );
  BUFX2 U10587 ( .A(n31314), .Y(n22440) );
  BUFX2 U10588 ( .A(n31332), .Y(n22443) );
  BUFX2 U10589 ( .A(n31352), .Y(n22446) );
  BUFX2 U10590 ( .A(n31372), .Y(n22449) );
  BUFX2 U10591 ( .A(n31392), .Y(n22452) );
  BUFX2 U10592 ( .A(n31604), .Y(n22455) );
  BUFX2 U10593 ( .A(n31623), .Y(n22458) );
  BUFX2 U10594 ( .A(n31641), .Y(n22461) );
  BUFX2 U10595 ( .A(n31659), .Y(n22464) );
  BUFX2 U10596 ( .A(n31666), .Y(n22467) );
  BUFX2 U10597 ( .A(n31697), .Y(n22470) );
  BUFX2 U10598 ( .A(n31704), .Y(n22473) );
  BUFX2 U10599 ( .A(n31737), .Y(n22476) );
  BUFX2 U10600 ( .A(n31775), .Y(n22479) );
  BUFX2 U10601 ( .A(n31782), .Y(n22482) );
  BUFX2 U10602 ( .A(n31814), .Y(n22485) );
  BUFX2 U10603 ( .A(n31821), .Y(n22488) );
  BUFX2 U10604 ( .A(n31854), .Y(n22491) );
  BUFX2 U10605 ( .A(n31898), .Y(n22494) );
  BUFX2 U10606 ( .A(n31906), .Y(n22497) );
  BUFX2 U10607 ( .A(n32483), .Y(n22500) );
  BUFX2 U10608 ( .A(n32494), .Y(n22503) );
  BUFX2 U10609 ( .A(n32532), .Y(n22506) );
  BUFX2 U10610 ( .A(n32625), .Y(n22509) );
  BUFX2 U10611 ( .A(n32642), .Y(n22512) );
  BUFX2 U10612 ( .A(n32673), .Y(n22515) );
  BUFX2 U10613 ( .A(n32720), .Y(n22518) );
  BUFX2 U10614 ( .A(n32767), .Y(n22521) );
  BUFX2 U10615 ( .A(n32817), .Y(n22524) );
  BUFX2 U10616 ( .A(n32907), .Y(n22527) );
  BUFX2 U10617 ( .A(n32983), .Y(n22530) );
  BUFX2 U10618 ( .A(n33437), .Y(n22533) );
  BUFX2 U10619 ( .A(n33440), .Y(n22536) );
  BUFX2 U10620 ( .A(n33443), .Y(n22539) );
  BUFX2 U10621 ( .A(n33455), .Y(n22542) );
  BUFX2 U10622 ( .A(n33458), .Y(n22545) );
  BUFX2 U10623 ( .A(n33461), .Y(n22548) );
  BUFX2 U10624 ( .A(n33465), .Y(n22551) );
  BUFX2 U10625 ( .A(n33501), .Y(n22554) );
  BUFX2 U10626 ( .A(n33504), .Y(n22557) );
  BUFX2 U10627 ( .A(n33507), .Y(n22560) );
  BUFX2 U10628 ( .A(n33534), .Y(n22563) );
  BUFX2 U10629 ( .A(n33541), .Y(n22566) );
  BUFX2 U10630 ( .A(n33547), .Y(n22569) );
  BUFX2 U10631 ( .A(n33550), .Y(n22572) );
  BUFX2 U10632 ( .A(n33554), .Y(n22575) );
  BUFX2 U10633 ( .A(n33580), .Y(n22578) );
  BUFX2 U10634 ( .A(n33583), .Y(n22581) );
  BUFX2 U10635 ( .A(n33586), .Y(n22584) );
  BUFX2 U10636 ( .A(n33590), .Y(n22587) );
  BUFX2 U10637 ( .A(n33602), .Y(n22590) );
  BUFX2 U10638 ( .A(n33605), .Y(n22593) );
  BUFX2 U10639 ( .A(n33608), .Y(n22596) );
  BUFX2 U10640 ( .A(n33612), .Y(n22599) );
  BUFX2 U10641 ( .A(n33624), .Y(n22602) );
  BUFX2 U10642 ( .A(n33627), .Y(n22605) );
  BUFX2 U10643 ( .A(n33630), .Y(n22608) );
  BUFX2 U10644 ( .A(n33633), .Y(n22611) );
  BUFX2 U10645 ( .A(n33646), .Y(n22614) );
  BUFX2 U10646 ( .A(n33649), .Y(n22617) );
  BUFX2 U10647 ( .A(n33652), .Y(n22620) );
  BUFX2 U10648 ( .A(n33656), .Y(n22623) );
  BUFX2 U10649 ( .A(n33668), .Y(n22638) );
  BUFX2 U10650 ( .A(n33671), .Y(n22639) );
  BUFX2 U10651 ( .A(n33674), .Y(n22640) );
  BUFX2 U10652 ( .A(n33689), .Y(n22641) );
  BUFX2 U10653 ( .A(n33695), .Y(n22642) );
  BUFX2 U10654 ( .A(n33711), .Y(n22643) );
  BUFX2 U10655 ( .A(n33717), .Y(n22644) );
  BUFX2 U10656 ( .A(n33733), .Y(n22645) );
  BUFX2 U10657 ( .A(n33739), .Y(n22646) );
  BUFX2 U10658 ( .A(n33755), .Y(n22647) );
  BUFX2 U10659 ( .A(n33761), .Y(n22648) );
  BUFX2 U10660 ( .A(n33777), .Y(n22649) );
  BUFX2 U10661 ( .A(n33783), .Y(n22650) );
  BUFX2 U10662 ( .A(n33915), .Y(n22651) );
  BUFX2 U10663 ( .A(n34195), .Y(n22652) );
  BUFX2 U10664 ( .A(n30898), .Y(n22653) );
  BUFX2 U10665 ( .A(n31465), .Y(n22654) );
  BUFX2 U10666 ( .A(n31920), .Y(n22655) );
  BUFX2 U10667 ( .A(n31932), .Y(n22656) );
  BUFX2 U10668 ( .A(n31942), .Y(n22657) );
  BUFX2 U10669 ( .A(n31952), .Y(n22658) );
  BUFX2 U10670 ( .A(n31963), .Y(n22659) );
  BUFX2 U10671 ( .A(n31973), .Y(n22660) );
  BUFX2 U10672 ( .A(n31982), .Y(n22661) );
  BUFX2 U10673 ( .A(n31993), .Y(n22662) );
  BUFX2 U10674 ( .A(n32049), .Y(n22663) );
  BUFX2 U10675 ( .A(n32057), .Y(n22664) );
  BUFX2 U10676 ( .A(n32064), .Y(n22665) );
  BUFX2 U10677 ( .A(n32072), .Y(n22666) );
  BUFX2 U10678 ( .A(n32080), .Y(n22667) );
  BUFX2 U10679 ( .A(n32088), .Y(n22668) );
  BUFX2 U10680 ( .A(n32095), .Y(n22669) );
  BUFX2 U10681 ( .A(n32105), .Y(n22670) );
  OR2X2 U10682 ( .A(n24015), .B(n25517), .Y(n32844) );
  INVX1 U10683 ( .A(n32844), .Y(n22671) );
  AND2X2 U10684 ( .A(n24977), .B(n23645), .Y(n34381) );
  INVX1 U10685 ( .A(n34381), .Y(n22672) );
  BUFX2 U10686 ( .A(n25716), .Y(n22673) );
  BUFX2 U10687 ( .A(n29485), .Y(n22674) );
  BUFX2 U10688 ( .A(n30137), .Y(n22675) );
  BUFX2 U10689 ( .A(n32801), .Y(n22676) );
  BUFX2 U10690 ( .A(n34255), .Y(n22677) );
  AND2X2 U10691 ( .A(n29590), .B(n29579), .Y(n33993) );
  AND2X2 U10692 ( .A(n29933), .B(n21106), .Y(n29836) );
  AND2X2 U10693 ( .A(n29902), .B(n25723), .Y(n32490) );
  BUFX2 U10694 ( .A(n33173), .Y(n22678) );
  AND2X2 U10695 ( .A(T[4]), .B(n34293), .Y(n25213) );
  INVX1 U10696 ( .A(n25213), .Y(n22679) );
  AND2X2 U10697 ( .A(net95147), .B(net104479), .Y(n33178) );
  INVX1 U10698 ( .A(n33178), .Y(n22680) );
  AND2X2 U10699 ( .A(n21219), .B(net149936), .Y(n33180) );
  INVX1 U10700 ( .A(n33180), .Y(n22681) );
  AND2X2 U10701 ( .A(net95147), .B(net124030), .Y(n33190) );
  INVX1 U10702 ( .A(n33190), .Y(n22682) );
  AND2X2 U10703 ( .A(net95147), .B(n28220), .Y(n33193) );
  INVX1 U10704 ( .A(n33193), .Y(n22683) );
  BUFX2 U10705 ( .A(n33070), .Y(n22684) );
  BUFX2 U10706 ( .A(n33083), .Y(n22685) );
  BUFX2 U10707 ( .A(n34176), .Y(n22686) );
  BUFX2 U10708 ( .A(n34297), .Y(n22687) );
  OR2X2 U10709 ( .A(n21187), .B(n21076), .Y(n29493) );
  INVX1 U10710 ( .A(n29493), .Y(n22688) );
  AND2X1 U10711 ( .A(n29387), .B(n26879), .Y(n33182) );
  INVX1 U10712 ( .A(n33182), .Y(n22689) );
  AND2X2 U10713 ( .A(n29416), .B(n21387), .Y(n33208) );
  INVX1 U10714 ( .A(n33208), .Y(n22690) );
  AND2X2 U10715 ( .A(n29391), .B(n21387), .Y(n33217) );
  INVX1 U10716 ( .A(n33217), .Y(n22691) );
  AND2X2 U10717 ( .A(n29415), .B(n33246), .Y(n33239) );
  INVX1 U10718 ( .A(n33239), .Y(n22692) );
  AND2X2 U10719 ( .A(n29391), .B(n33246), .Y(n33248) );
  INVX1 U10720 ( .A(n33248), .Y(n22693) );
  AND2X2 U10721 ( .A(n29415), .B(n25430), .Y(n33269) );
  INVX1 U10722 ( .A(n33269), .Y(n22694) );
  AND2X2 U10723 ( .A(n29391), .B(n25430), .Y(n33278) );
  INVX1 U10724 ( .A(n33278), .Y(n22695) );
  AND2X2 U10725 ( .A(n29415), .B(n25429), .Y(n33300) );
  INVX1 U10726 ( .A(n33300), .Y(n22696) );
  AND2X2 U10727 ( .A(n29391), .B(n25429), .Y(n33309) );
  INVX1 U10728 ( .A(n33309), .Y(n22697) );
  AND2X2 U10729 ( .A(n29415), .B(n33338), .Y(n33331) );
  INVX1 U10730 ( .A(n33331), .Y(n22698) );
  AND2X2 U10731 ( .A(n29391), .B(n33338), .Y(n33340) );
  INVX1 U10732 ( .A(n33340), .Y(n22699) );
  AND2X2 U10733 ( .A(n29415), .B(n33368), .Y(n33361) );
  INVX1 U10734 ( .A(n33361), .Y(n22700) );
  AND2X1 U10735 ( .A(n29391), .B(n33368), .Y(n33370) );
  INVX1 U10736 ( .A(n33370), .Y(n22701) );
  AND2X2 U10737 ( .A(n29415), .B(n21384), .Y(n33391) );
  INVX1 U10738 ( .A(n33391), .Y(n22702) );
  AND2X2 U10739 ( .A(n29391), .B(n21384), .Y(n33400) );
  INVX1 U10740 ( .A(n33400), .Y(n22703) );
  AND2X2 U10741 ( .A(n29415), .B(n25773), .Y(n33422) );
  INVX1 U10742 ( .A(n33422), .Y(n22704) );
  AND2X2 U10743 ( .A(n29391), .B(n25773), .Y(n33431) );
  INVX1 U10744 ( .A(n33431), .Y(n22705) );
  AND2X2 U10745 ( .A(n29415), .B(n25427), .Y(n33466) );
  INVX1 U10746 ( .A(n33466), .Y(n22706) );
  AND2X2 U10747 ( .A(n29415), .B(n25456), .Y(n33512) );
  INVX1 U10748 ( .A(n33512), .Y(n22707) );
  AND2X2 U10749 ( .A(n29415), .B(n25424), .Y(n33568) );
  INVX1 U10750 ( .A(n33568), .Y(n22708) );
  AND2X2 U10751 ( .A(n29415), .B(n25432), .Y(n33591) );
  INVX1 U10752 ( .A(n33591), .Y(n22709) );
  AND2X2 U10753 ( .A(n29415), .B(n26940), .Y(n33613) );
  INVX1 U10754 ( .A(n33613), .Y(n22710) );
  AND2X2 U10755 ( .A(n29415), .B(n25440), .Y(n33634) );
  INVX1 U10756 ( .A(n33634), .Y(n22711) );
  AND2X2 U10757 ( .A(n29416), .B(n33682), .Y(n33678) );
  INVX1 U10758 ( .A(n33678), .Y(n22712) );
  AND2X2 U10759 ( .A(n29416), .B(n26942), .Y(n33700) );
  INVX1 U10760 ( .A(n33700), .Y(n22713) );
  AND2X2 U10761 ( .A(n29415), .B(n26765), .Y(n33722) );
  INVX1 U10762 ( .A(n33722), .Y(n22714) );
  AND2X2 U10763 ( .A(n29415), .B(n23111), .Y(n33743) );
  INVX1 U10764 ( .A(n33743), .Y(n22715) );
  AND2X2 U10765 ( .A(n29416), .B(n27021), .Y(n33810) );
  INVX1 U10766 ( .A(n33810), .Y(n22716) );
  AND2X2 U10767 ( .A(n29416), .B(n26820), .Y(n33879) );
  INVX1 U10768 ( .A(n33879), .Y(n22717) );
  AND2X2 U10769 ( .A(n29387), .B(n26820), .Y(n33886) );
  INVX1 U10770 ( .A(n33886), .Y(n22718) );
  OR2X2 U10771 ( .A(n25615), .B(n34196), .Y(n33926) );
  INVX1 U10772 ( .A(n33926), .Y(n22719) );
  AND2X2 U10773 ( .A(n29417), .B(n26879), .Y(n34220) );
  INVX1 U10774 ( .A(n34220), .Y(n22720) );
  OR2X2 U10775 ( .A(n21105), .B(n34310), .Y(n34300) );
  INVX1 U10776 ( .A(n34300), .Y(n22721) );
  BUFX2 U10777 ( .A(n33150), .Y(n22722) );
  AND2X2 U10778 ( .A(n21420), .B(n21551), .Y(n34188) );
  INVX1 U10779 ( .A(n34188), .Y(n22723) );
  AND2X2 U10780 ( .A(n21537), .B(n34180), .Y(n34182) );
  INVX1 U10781 ( .A(n34182), .Y(n22724) );
  BUFX2 U10782 ( .A(n33101), .Y(n22725) );
  AND2X2 U10783 ( .A(n23103), .B(n23200), .Y(n29585) );
  INVX1 U10784 ( .A(n29585), .Y(n22726) );
  BUFX2 U10785 ( .A(n30669), .Y(n22727) );
  OR2X2 U10786 ( .A(n22109), .B(n22129), .Y(n29538) );
  INVX1 U10787 ( .A(n29538), .Y(n22728) );
  AND2X2 U10788 ( .A(n25915), .B(n32434), .Y(n31760) );
  INVX1 U10789 ( .A(n31760), .Y(n22729) );
  INVX1 U10790 ( .A(n32198), .Y(n22730) );
  AND2X2 U10791 ( .A(n3275), .B(n32764), .Y(n32766) );
  INVX1 U10792 ( .A(n32766), .Y(n22731) );
  AND2X2 U10793 ( .A(n3151), .B(n21212), .Y(n32984) );
  INVX1 U10794 ( .A(n32984), .Y(n22732) );
  AND2X2 U10795 ( .A(n20956), .B(n27178), .Y(n34294) );
  INVX1 U10796 ( .A(n34294), .Y(n22733) );
  BUFX2 U10797 ( .A(n29599), .Y(n22734) );
  BUFX2 U10798 ( .A(n30662), .Y(n22735) );
  BUFX2 U10799 ( .A(n30705), .Y(n22736) );
  BUFX2 U10800 ( .A(n30725), .Y(n22737) );
  BUFX2 U10801 ( .A(n30744), .Y(n22738) );
  BUFX2 U10802 ( .A(n30765), .Y(n22739) );
  BUFX2 U10803 ( .A(n30784), .Y(n22740) );
  BUFX2 U10804 ( .A(n30805), .Y(n22741) );
  BUFX2 U10805 ( .A(n30824), .Y(n22742) );
  BUFX2 U10806 ( .A(n31218), .Y(n22743) );
  BUFX2 U10807 ( .A(n31258), .Y(n22744) );
  BUFX2 U10808 ( .A(n31412), .Y(n22745) );
  BUFX2 U10809 ( .A(n31433), .Y(n22746) );
  BUFX2 U10810 ( .A(n31452), .Y(n22747) );
  BUFX2 U10811 ( .A(n32492), .Y(n22748) );
  BUFX2 U10812 ( .A(n32550), .Y(n22749) );
  BUFX2 U10813 ( .A(n32765), .Y(n22750) );
  BUFX2 U10814 ( .A(n32917), .Y(n22751) );
  BUFX2 U10815 ( .A(n32985), .Y(n22752) );
  BUFX2 U10816 ( .A(n33478), .Y(n22753) );
  BUFX2 U10817 ( .A(n33481), .Y(n22754) );
  BUFX2 U10818 ( .A(n33484), .Y(n22755) );
  BUFX2 U10819 ( .A(n33488), .Y(n22756) );
  BUFX2 U10820 ( .A(n33511), .Y(n22757) );
  BUFX2 U10821 ( .A(n33524), .Y(n22758) );
  BUFX2 U10822 ( .A(n33527), .Y(n22759) );
  BUFX2 U10823 ( .A(n33530), .Y(n22760) );
  BUFX2 U10824 ( .A(n33537), .Y(n22761) );
  BUFX2 U10825 ( .A(n33544), .Y(n22762) );
  BUFX2 U10826 ( .A(n33675), .Y(n22763) );
  BUFX2 U10827 ( .A(n33690), .Y(n22764) );
  BUFX2 U10828 ( .A(n33697), .Y(n22765) );
  BUFX2 U10829 ( .A(n33712), .Y(n22766) );
  BUFX2 U10830 ( .A(n33719), .Y(n22767) );
  BUFX2 U10831 ( .A(n33734), .Y(n22768) );
  BUFX2 U10832 ( .A(n33740), .Y(n22769) );
  BUFX2 U10833 ( .A(n33756), .Y(n22770) );
  BUFX2 U10834 ( .A(n33763), .Y(n22771) );
  BUFX2 U10835 ( .A(n33778), .Y(n22772) );
  BUFX2 U10836 ( .A(n33785), .Y(n22773) );
  BUFX2 U10837 ( .A(n33797), .Y(n22774) );
  BUFX2 U10838 ( .A(n33800), .Y(n22775) );
  BUFX2 U10839 ( .A(n33803), .Y(n22776) );
  BUFX2 U10840 ( .A(n33807), .Y(n22777) );
  BUFX2 U10841 ( .A(n33820), .Y(n22778) );
  BUFX2 U10842 ( .A(n33823), .Y(n22779) );
  BUFX2 U10843 ( .A(n33826), .Y(n22780) );
  BUFX2 U10844 ( .A(n33830), .Y(n22781) );
  BUFX2 U10845 ( .A(n33843), .Y(n22782) );
  BUFX2 U10846 ( .A(n33846), .Y(n22783) );
  BUFX2 U10847 ( .A(n33849), .Y(n22784) );
  BUFX2 U10848 ( .A(n33853), .Y(n22785) );
  BUFX2 U10849 ( .A(n33866), .Y(n22786) );
  BUFX2 U10850 ( .A(n33869), .Y(n22787) );
  BUFX2 U10851 ( .A(n33872), .Y(n22788) );
  BUFX2 U10852 ( .A(n33876), .Y(n22789) );
  BUFX2 U10853 ( .A(n33891), .Y(n22790) );
  BUFX2 U10854 ( .A(n33894), .Y(n22791) );
  BUFX2 U10855 ( .A(n33897), .Y(n22792) );
  BUFX2 U10856 ( .A(n33901), .Y(n22793) );
  BUFX2 U10857 ( .A(n31913), .Y(n22794) );
  BUFX2 U10858 ( .A(n30647), .Y(n22795) );
  BUFX2 U10859 ( .A(n30838), .Y(n22796) );
  BUFX2 U10860 ( .A(n30878), .Y(n22797) );
  BUFX2 U10861 ( .A(n30959), .Y(n22798) );
  BUFX2 U10862 ( .A(n31054), .Y(n22799) );
  BUFX2 U10863 ( .A(n31134), .Y(n22800) );
  BUFX2 U10864 ( .A(n31172), .Y(n22801) );
  BUFX2 U10865 ( .A(n31289), .Y(n22802) );
  BUFX2 U10866 ( .A(n31308), .Y(n22803) );
  BUFX2 U10867 ( .A(n31325), .Y(n22804) );
  BUFX2 U10868 ( .A(n31345), .Y(n22805) );
  BUFX2 U10869 ( .A(n31365), .Y(n22806) );
  BUFX2 U10870 ( .A(n31385), .Y(n22807) );
  BUFX2 U10871 ( .A(n31405), .Y(n22808) );
  BUFX2 U10872 ( .A(n31426), .Y(n22809) );
  BUFX2 U10873 ( .A(n31446), .Y(n22810) );
  BUFX2 U10874 ( .A(n31485), .Y(n22811) );
  BUFX2 U10875 ( .A(n31522), .Y(n22812) );
  BUFX2 U10876 ( .A(n31754), .Y(n22813) );
  BUFX2 U10877 ( .A(n31794), .Y(n22814) );
  BUFX2 U10878 ( .A(n31833), .Y(n22815) );
  BUFX2 U10879 ( .A(n31873), .Y(n22816) );
  OR2X2 U10880 ( .A(n23473), .B(n23474), .Y(n33025) );
  OR2X2 U10881 ( .A(n30690), .B(n30689), .Y(n30691) );
  INVX1 U10882 ( .A(n30691), .Y(n22817) );
  OR2X2 U10883 ( .A(n30707), .B(n30709), .Y(n30710) );
  INVX1 U10884 ( .A(n30710), .Y(n22818) );
  OR2X2 U10885 ( .A(n30727), .B(n30729), .Y(n30730) );
  INVX1 U10886 ( .A(n30730), .Y(n22819) );
  OR2X2 U10887 ( .A(n30749), .B(n30748), .Y(n30750) );
  INVX1 U10888 ( .A(n30750), .Y(n22820) );
  OR2X2 U10889 ( .A(n30767), .B(n30769), .Y(n30770) );
  INVX1 U10890 ( .A(n30770), .Y(n22821) );
  OR2X2 U10891 ( .A(n30789), .B(n30788), .Y(n30790) );
  INVX1 U10892 ( .A(n30790), .Y(n22822) );
  OR2X2 U10893 ( .A(n30807), .B(n30809), .Y(n30810) );
  INVX1 U10894 ( .A(n30810), .Y(n22823) );
  OR2X2 U10895 ( .A(n30829), .B(n30828), .Y(n30830) );
  INVX1 U10896 ( .A(n30830), .Y(n22824) );
  OR2X2 U10897 ( .A(n30847), .B(n30849), .Y(n30850) );
  INVX1 U10898 ( .A(n30850), .Y(n22825) );
  OR2X2 U10899 ( .A(n30869), .B(n30868), .Y(n30870) );
  INVX1 U10900 ( .A(n30870), .Y(n22826) );
  OR2X2 U10901 ( .A(n30890), .B(n30889), .Y(n30891) );
  INVX1 U10902 ( .A(n30891), .Y(n22827) );
  OR2X2 U10903 ( .A(n30910), .B(n30909), .Y(n30911) );
  INVX1 U10904 ( .A(n30911), .Y(n22828) );
  OR2X2 U10905 ( .A(n30928), .B(n30930), .Y(n30931) );
  INVX1 U10906 ( .A(n30931), .Y(n22829) );
  OR2X2 U10907 ( .A(n30950), .B(n30949), .Y(n30951) );
  INVX1 U10908 ( .A(n30951), .Y(n22830) );
  OR2X2 U10909 ( .A(n30971), .B(n30970), .Y(n30972) );
  INVX1 U10910 ( .A(n30972), .Y(n22831) );
  OR2X2 U10911 ( .A(n30991), .B(n30990), .Y(n30992) );
  INVX1 U10912 ( .A(n30992), .Y(n22832) );
  OR2X2 U10913 ( .A(n27230), .B(n31007), .Y(n31008) );
  INVX1 U10914 ( .A(n31008), .Y(n22833) );
  OR2X2 U10915 ( .A(n31028), .B(n31027), .Y(n31029) );
  INVX1 U10916 ( .A(n31029), .Y(n22834) );
  OR2X2 U10917 ( .A(n27231), .B(n31045), .Y(n31046) );
  INVX1 U10918 ( .A(n31046), .Y(n22835) );
  OR2X2 U10919 ( .A(n31066), .B(n31065), .Y(n31067) );
  INVX1 U10920 ( .A(n31067), .Y(n22836) );
  OR2X2 U10921 ( .A(n31085), .B(n31084), .Y(n31086) );
  INVX1 U10922 ( .A(n31086), .Y(n22837) );
  OR2X2 U10923 ( .A(n31106), .B(n31105), .Y(n31107) );
  INVX1 U10924 ( .A(n31107), .Y(n22838) );
  OR2X2 U10925 ( .A(n31125), .B(n31124), .Y(n31126) );
  INVX1 U10926 ( .A(n31126), .Y(n22839) );
  OR2X2 U10927 ( .A(n31146), .B(n31145), .Y(n31147) );
  INVX1 U10928 ( .A(n31147), .Y(n22840) );
  OR2X2 U10929 ( .A(n27228), .B(n31163), .Y(n31164) );
  INVX1 U10930 ( .A(n31164), .Y(n22841) );
  OR2X2 U10931 ( .A(n31183), .B(n31182), .Y(n31184) );
  INVX1 U10932 ( .A(n31184), .Y(n22842) );
  OR2X2 U10933 ( .A(n31202), .B(n31201), .Y(n31203) );
  INVX1 U10934 ( .A(n31203), .Y(n22843) );
  OR2X2 U10935 ( .A(n31222), .B(n31223), .Y(n31224) );
  INVX1 U10936 ( .A(n31224), .Y(n22844) );
  OR2X2 U10937 ( .A(n31242), .B(n31241), .Y(n31243) );
  INVX1 U10938 ( .A(n31243), .Y(n22845) );
  OR2X2 U10939 ( .A(n31263), .B(n31262), .Y(n31264) );
  INVX1 U10940 ( .A(n31264), .Y(n22846) );
  OR2X2 U10941 ( .A(n31274), .B(n31281), .Y(n31282) );
  INVX1 U10942 ( .A(n31282), .Y(n22847) );
  OR2X2 U10943 ( .A(n31297), .B(n31299), .Y(n31300) );
  INVX1 U10944 ( .A(n31300), .Y(n22848) );
  OR2X2 U10945 ( .A(n31316), .B(n31317), .Y(n31318) );
  INVX1 U10946 ( .A(n31318), .Y(n22849) );
  OR2X2 U10947 ( .A(n31334), .B(n31336), .Y(n31337) );
  INVX1 U10948 ( .A(n31337), .Y(n22850) );
  OR2X2 U10949 ( .A(n31357), .B(n31356), .Y(n31358) );
  INVX1 U10950 ( .A(n31358), .Y(n22851) );
  OR2X2 U10951 ( .A(n31374), .B(n31376), .Y(n31377) );
  INVX1 U10952 ( .A(n31377), .Y(n22852) );
  OR2X2 U10953 ( .A(n31396), .B(n31397), .Y(n31398) );
  INVX1 U10954 ( .A(n31398), .Y(n22853) );
  OR2X2 U10955 ( .A(n31417), .B(n31416), .Y(n31418) );
  INVX1 U10956 ( .A(n31418), .Y(n22854) );
  OR2X2 U10957 ( .A(n31438), .B(n31437), .Y(n31439) );
  INVX1 U10958 ( .A(n31439), .Y(n22855) );
  OR2X2 U10959 ( .A(n31454), .B(n31456), .Y(n31457) );
  INVX1 U10960 ( .A(n31457), .Y(n22856) );
  OR2X2 U10961 ( .A(n31477), .B(n31476), .Y(n31478) );
  INVX1 U10962 ( .A(n31478), .Y(n22857) );
  OR2X2 U10963 ( .A(n31494), .B(n31495), .Y(n31496) );
  INVX1 U10964 ( .A(n31496), .Y(n22858) );
  OR2X2 U10965 ( .A(n25460), .B(n31514), .Y(n31515) );
  INVX1 U10966 ( .A(n31515), .Y(n22859) );
  OR2X2 U10967 ( .A(n31531), .B(n31533), .Y(n31534) );
  INVX1 U10968 ( .A(n31534), .Y(n22860) );
  OR2X2 U10969 ( .A(n31554), .B(n31553), .Y(n31555) );
  INVX1 U10970 ( .A(n31555), .Y(n22861) );
  OR2X2 U10971 ( .A(n31574), .B(n31573), .Y(n31575) );
  INVX1 U10972 ( .A(n31575), .Y(n22862) );
  OR2X2 U10973 ( .A(n31592), .B(n31594), .Y(n31595) );
  INVX1 U10974 ( .A(n31595), .Y(n22863) );
  OR2X2 U10975 ( .A(n31614), .B(n31613), .Y(n31615) );
  INVX1 U10976 ( .A(n31615), .Y(n22864) );
  OR2X2 U10977 ( .A(n27226), .B(n31631), .Y(n31632) );
  INVX1 U10978 ( .A(n31632), .Y(n22865) );
  INVX1 U10979 ( .A(n31651), .Y(n22866) );
  INVX1 U10980 ( .A(n31669), .Y(n22867) );
  OR2X2 U10981 ( .A(n31686), .B(n31688), .Y(n31689) );
  INVX1 U10982 ( .A(n31689), .Y(n22868) );
  OR2X2 U10983 ( .A(n31707), .B(n31706), .Y(n31708) );
  INVX1 U10984 ( .A(n31708), .Y(n22869) );
  OR2X2 U10985 ( .A(n31728), .B(n31727), .Y(n31729) );
  INVX1 U10986 ( .A(n31729), .Y(n22870) );
  OR2X2 U10987 ( .A(n27227), .B(n31745), .Y(n31746) );
  INVX1 U10988 ( .A(n31746), .Y(n22871) );
  OR2X2 U10989 ( .A(n31766), .B(n31765), .Y(n31767) );
  INVX1 U10990 ( .A(n31767), .Y(n22872) );
  OR2X2 U10991 ( .A(n31785), .B(n31784), .Y(n31786) );
  INVX1 U10992 ( .A(n31786), .Y(n22873) );
  OR2X2 U10993 ( .A(n31803), .B(n31805), .Y(n31806) );
  INVX1 U10994 ( .A(n31806), .Y(n22874) );
  OR2X2 U10995 ( .A(n31824), .B(n31823), .Y(n31825) );
  INVX1 U10996 ( .A(n31825), .Y(n22875) );
  OR2X2 U10997 ( .A(n31842), .B(n31844), .Y(n31845) );
  INVX1 U10998 ( .A(n31845), .Y(n22876) );
  OR2X2 U10999 ( .A(n27229), .B(n31863), .Y(n31864) );
  INVX1 U11000 ( .A(n31864), .Y(n22877) );
  OR2X2 U11001 ( .A(n31883), .B(n31886), .Y(n31887) );
  INVX1 U11002 ( .A(n31887), .Y(n22878) );
  AND2X2 U11003 ( .A(n25206), .B(n25196), .Y(n33124) );
  INVX1 U11004 ( .A(n33124), .Y(n22879) );
  AND2X2 U11005 ( .A(n34330), .B(n34407), .Y(n34327) );
  AND2X2 U11006 ( .A(n34435), .B(n34434), .Y(n34436) );
  AND2X2 U11007 ( .A(n29484), .B(n21067), .Y(n7906) );
  INVX1 U11008 ( .A(n7906), .Y(n22880) );
  INVX1 U11009 ( .A(n7906), .Y(n22881) );
  BUFX2 U11010 ( .A(n32488), .Y(n22882) );
  INVX1 U11011 ( .A(n32502), .Y(n22884) );
  INVX1 U11012 ( .A(n32504), .Y(n22885) );
  BUFX2 U11013 ( .A(n32540), .Y(n22887) );
  BUFX2 U11014 ( .A(n32559), .Y(n22888) );
  INVX1 U11015 ( .A(n32578), .Y(n22890) );
  INVX1 U11016 ( .A(n32580), .Y(n22891) );
  INVX1 U11017 ( .A(n32600), .Y(n22894) );
  BUFX2 U11018 ( .A(n32680), .Y(n22896) );
  INVX1 U11019 ( .A(n32681), .Y(n22898) );
  INVX1 U11020 ( .A(n32683), .Y(n22899) );
  INVX1 U11021 ( .A(n32690), .Y(n22902) );
  INVX1 U11022 ( .A(n32692), .Y(n22903) );
  BUFX2 U11023 ( .A(n32727), .Y(n22905) );
  INVX1 U11024 ( .A(n32787), .Y(n22907) );
  INVX1 U11025 ( .A(n32789), .Y(n22908) );
  INVX1 U11026 ( .A(n32859), .Y(n22911) );
  INVX1 U11027 ( .A(n32861), .Y(n22912) );
  INVX1 U11028 ( .A(n32867), .Y(n22915) );
  INVX1 U11029 ( .A(n32869), .Y(n22916) );
  BUFX2 U11030 ( .A(n32916), .Y(n22918) );
  BUFX2 U11031 ( .A(n32925), .Y(n22919) );
  INVX1 U11032 ( .A(n32958), .Y(n22921) );
  INVX1 U11033 ( .A(n32960), .Y(n22922) );
  INVX1 U11034 ( .A(n32974), .Y(n22925) );
  INVX1 U11035 ( .A(n32975), .Y(n22926) );
  BUFX2 U11036 ( .A(n33024), .Y(n22927) );
  AND2X2 U11037 ( .A(n21528), .B(n24880), .Y(n32549) );
  INVX1 U11038 ( .A(n32549), .Y(n22928) );
  INVX1 U11039 ( .A(n32641), .Y(n22929) );
  AND2X2 U11040 ( .A(n21530), .B(n24884), .Y(n32831) );
  INVX1 U11041 ( .A(n32831), .Y(n22930) );
  AND2X2 U11042 ( .A(n21531), .B(n24885), .Y(n32934) );
  INVX1 U11043 ( .A(n32934), .Y(n22931) );
  AND2X2 U11044 ( .A(n21532), .B(n24886), .Y(n33043) );
  INVX1 U11045 ( .A(n33043), .Y(n22932) );
  AND2X2 U11046 ( .A(n29510), .B(n25763), .Y(n29505) );
  INVX1 U11047 ( .A(n29505), .Y(n22933) );
  INVX1 U11048 ( .A(n32778), .Y(n22935) );
  INVX1 U11049 ( .A(n32780), .Y(n22936) );
  AND2X2 U11050 ( .A(n25714), .B(n34441), .Y(n25733) );
  INVX1 U11051 ( .A(n25733), .Y(n22938) );
  AND2X2 U11052 ( .A(n27117), .B(n29526), .Y(n34613) );
  INVX1 U11053 ( .A(n34613), .Y(n22939) );
  AND2X2 U11054 ( .A(n23283), .B(n21106), .Y(n33904) );
  INVX1 U11055 ( .A(n33904), .Y(n22940) );
  INVX1 U11056 ( .A(n33904), .Y(n22941) );
  AND2X2 U11057 ( .A(n22941), .B(n26820), .Y(n33890) );
  INVX1 U11058 ( .A(n33890), .Y(n22942) );
  AND2X2 U11059 ( .A(n23111), .B(n25770), .Y(n30514) );
  INVX1 U11060 ( .A(n30514), .Y(n22943) );
  AND2X2 U11061 ( .A(n26765), .B(n27027), .Y(n30519) );
  INVX1 U11062 ( .A(n30519), .Y(n22944) );
  AND2X2 U11063 ( .A(n25440), .B(n32953), .Y(n30536) );
  INVX1 U11064 ( .A(n30536), .Y(n22945) );
  AND2X2 U11065 ( .A(n26940), .B(n27024), .Y(n30541) );
  INVX1 U11066 ( .A(n30541), .Y(n22946) );
  AND2X2 U11067 ( .A(n23446), .B(n21106), .Y(n29871) );
  INVX1 U11068 ( .A(n29871), .Y(n22947) );
  INVX1 U11069 ( .A(n29871), .Y(n22948) );
  AND2X2 U11070 ( .A(n25432), .B(n22948), .Y(n30546) );
  INVX1 U11071 ( .A(n30546), .Y(n22949) );
  AND2X2 U11072 ( .A(n25403), .B(n25597), .Y(n29886) );
  INVX1 U11073 ( .A(n29886), .Y(n22950) );
  AND2X2 U11074 ( .A(n25456), .B(n25202), .Y(n30558) );
  INVX1 U11075 ( .A(n30558), .Y(n22951) );
  AND2X2 U11076 ( .A(n25427), .B(n25351), .Y(n30567) );
  INVX1 U11077 ( .A(n30567), .Y(n22952) );
  AND2X2 U11078 ( .A(n25438), .B(n25347), .Y(n30572) );
  INVX1 U11079 ( .A(n30572), .Y(n22953) );
  AND2X2 U11080 ( .A(n25773), .B(n25350), .Y(n30577) );
  INVX1 U11081 ( .A(n30577), .Y(n22954) );
  AND2X2 U11082 ( .A(n21384), .B(n25353), .Y(n30582) );
  INVX1 U11083 ( .A(n30582), .Y(n22955) );
  AND2X2 U11084 ( .A(n33368), .B(n21435), .Y(n30587) );
  INVX1 U11085 ( .A(n30587), .Y(n22956) );
  AND2X2 U11086 ( .A(n33338), .B(n25453), .Y(n30592) );
  INVX1 U11087 ( .A(n30592), .Y(n22957) );
  AND2X2 U11088 ( .A(n25429), .B(n25355), .Y(n30597) );
  INVX1 U11089 ( .A(n30597), .Y(n22958) );
  AND2X2 U11090 ( .A(n25430), .B(n25442), .Y(n30602) );
  INVX1 U11091 ( .A(n30602), .Y(n22959) );
  AND2X2 U11092 ( .A(n33246), .B(n26269), .Y(n30607) );
  INVX1 U11093 ( .A(n30607), .Y(n22960) );
  AND2X2 U11094 ( .A(n21387), .B(n23112), .Y(n30612) );
  INVX1 U11095 ( .A(n30612), .Y(n22961) );
  BUFX2 U11096 ( .A(n25755), .Y(n22962) );
  BUFX2 U11097 ( .A(n2247), .Y(n22964) );
  BUFX2 U11098 ( .A(n30630), .Y(n22965) );
  BUFX2 U11099 ( .A(n32940), .Y(n22966) );
  BUFX2 U11100 ( .A(n33075), .Y(n22967) );
  AND2X2 U11101 ( .A(n21069), .B(n21012), .Y(n29489) );
  INVX1 U11102 ( .A(n30474), .Y(n22968) );
  AND2X2 U11103 ( .A(n29825), .B(n27315), .Y(n29990) );
  INVX1 U11104 ( .A(n29990), .Y(n22969) );
  AND2X2 U11105 ( .A(n29922), .B(n21106), .Y(n29824) );
  INVX1 U11106 ( .A(n29824), .Y(n22970) );
  AND2X2 U11107 ( .A(n31868), .B(n25765), .Y(n31894) );
  INVX1 U11108 ( .A(n31894), .Y(n22971) );
  AND2X2 U11109 ( .A(n33052), .B(n33051), .Y(n34443) );
  AND2X2 U11110 ( .A(n34356), .B(n33078), .Y(n33096) );
  AND2X2 U11111 ( .A(n23070), .B(n25446), .Y(n34265) );
  INVX1 U11112 ( .A(n34265), .Y(n22972) );
  INVX1 U11113 ( .A(n34265), .Y(n22973) );
  AND2X2 U11114 ( .A(n34425), .B(n25748), .Y(n34431) );
  INVX1 U11115 ( .A(n34431), .Y(n22974) );
  INVX1 U11116 ( .A(n32878), .Y(n22976) );
  INVX1 U11117 ( .A(n32880), .Y(n22977) );
  INVX1 U11118 ( .A(n25848), .Y(n22979) );
  BUFX2 U11119 ( .A(n15179), .Y(n22980) );
  INVX1 U11120 ( .A(n25843), .Y(n22981) );
  INVX1 U11121 ( .A(n25843), .Y(n22982) );
  BUFX2 U11122 ( .A(n34179), .Y(n22983) );
  AND2X2 U11123 ( .A(locTrig[2]), .B(n29484), .Y(n30684) );
  INVX1 U11124 ( .A(n30684), .Y(n22984) );
  INVX1 U11125 ( .A(n30684), .Y(n22985) );
  AND2X2 U11126 ( .A(n23282), .B(n21106), .Y(n34192) );
  INVX1 U11127 ( .A(n34192), .Y(n22986) );
  AND2X2 U11128 ( .A(n29376), .B(n21558), .Y(n31902) );
  INVX1 U11129 ( .A(n31902), .Y(n22987) );
  AND2X1 U11130 ( .A(n34386), .B(n34385), .Y(n25166) );
  INVX1 U11131 ( .A(n25166), .Y(n22988) );
  AND2X2 U11132 ( .A(net95105), .B(net109585), .Y(n30075) );
  INVX1 U11133 ( .A(n30075), .Y(n22989) );
  INVX1 U11134 ( .A(n30075), .Y(n22990) );
  AND2X2 U11135 ( .A(T[4]), .B(n34442), .Y(n33136) );
  INVX1 U11136 ( .A(n33136), .Y(n22991) );
  AND2X2 U11137 ( .A(n34357), .B(n34356), .Y(n34364) );
  INVX1 U11138 ( .A(n34364), .Y(n22992) );
  INVX1 U11139 ( .A(n34364), .Y(n22993) );
  BUFX2 U11140 ( .A(n14358), .Y(net143010) );
  BUFX2 U11141 ( .A(n15184), .Y(n22994) );
  BUFX2 U11142 ( .A(n34178), .Y(n22995) );
  AND2X2 U11143 ( .A(n26986), .B(n23278), .Y(n25343) );
  INVX1 U11144 ( .A(n25343), .Y(n22996) );
  INVX1 U11145 ( .A(n34373), .Y(n22997) );
  AND2X1 U11146 ( .A(n30645), .B(net96340), .Y(n30668) );
  INVX1 U11147 ( .A(n30668), .Y(n22998) );
  AND2X1 U11148 ( .A(n31714), .B(net96340), .Y(n31725) );
  INVX1 U11149 ( .A(n31725), .Y(n22999) );
  AND2X1 U11150 ( .A(n20953), .B(n34351), .Y(n34251) );
  INVX1 U11151 ( .A(n34251), .Y(n23000) );
  INVX1 U11152 ( .A(n34311), .Y(n23001) );
  INVX1 U11153 ( .A(n20828), .Y(n23002) );
  AND2X1 U11154 ( .A(n30735), .B(net96340), .Y(n30746) );
  INVX1 U11155 ( .A(n30746), .Y(n23003) );
  AND2X1 U11156 ( .A(n30756), .B(net96340), .Y(n30767) );
  INVX1 U11157 ( .A(n30767), .Y(n23004) );
  AND2X1 U11158 ( .A(n30775), .B(net96340), .Y(n30786) );
  INVX1 U11159 ( .A(n30786), .Y(n23005) );
  AND2X1 U11160 ( .A(n30796), .B(net96340), .Y(n30807) );
  INVX1 U11161 ( .A(n30807), .Y(n23006) );
  AND2X1 U11162 ( .A(n30815), .B(net96340), .Y(n30826) );
  INVX1 U11163 ( .A(n30826), .Y(n23007) );
  AND2X1 U11164 ( .A(n30836), .B(net96340), .Y(n30847) );
  INVX1 U11165 ( .A(n30847), .Y(n23008) );
  AND2X1 U11166 ( .A(n30876), .B(net96340), .Y(n30887) );
  INVX1 U11167 ( .A(n30887), .Y(n23009) );
  AND2X1 U11168 ( .A(n30896), .B(net96340), .Y(n30907) );
  INVX1 U11169 ( .A(n30907), .Y(n23010) );
  AND2X1 U11170 ( .A(n30936), .B(net96340), .Y(n30947) );
  INVX1 U11171 ( .A(n30947), .Y(n23012) );
  AND2X1 U11172 ( .A(n30957), .B(net96340), .Y(n30968) );
  INVX1 U11173 ( .A(n30968), .Y(n23013) );
  AND2X1 U11174 ( .A(n30978), .B(net96340), .Y(n30988) );
  INVX1 U11175 ( .A(n30988), .Y(n23014) );
  AND2X2 U11176 ( .A(n29376), .B(n30997), .Y(n31006) );
  INVX1 U11177 ( .A(n31006), .Y(n23015) );
  AND2X2 U11178 ( .A(n29376), .B(n31034), .Y(n31044) );
  INVX1 U11179 ( .A(n31044), .Y(n23016) );
  INVX1 U11180 ( .A(n31044), .Y(n23017) );
  AND2X1 U11181 ( .A(n31052), .B(net96340), .Y(n31063) );
  INVX1 U11182 ( .A(n31063), .Y(n23018) );
  AND2X2 U11183 ( .A(n29376), .B(n31072), .Y(n31083) );
  INVX1 U11184 ( .A(n31083), .Y(n23019) );
  AND2X1 U11185 ( .A(n31110), .B(net96340), .Y(n31117) );
  INVX1 U11186 ( .A(n31117), .Y(n23020) );
  AND2X2 U11187 ( .A(n25466), .B(n31112), .Y(n31123) );
  INVX1 U11188 ( .A(n31123), .Y(n23021) );
  INVX1 U11189 ( .A(n31123), .Y(n23022) );
  AND2X1 U11190 ( .A(n31132), .B(net96340), .Y(n31143) );
  INVX1 U11191 ( .A(n31143), .Y(n23023) );
  AND2X2 U11192 ( .A(n25466), .B(n21554), .Y(n31162) );
  INVX1 U11193 ( .A(n31162), .Y(n23024) );
  AND2X1 U11194 ( .A(n31170), .B(net96340), .Y(n31180) );
  INVX1 U11195 ( .A(n31180), .Y(n23025) );
  AND2X2 U11196 ( .A(n25466), .B(n31189), .Y(n31200) );
  INVX1 U11197 ( .A(n31200), .Y(n23026) );
  INVX1 U11198 ( .A(n31200), .Y(n23027) );
  AND2X1 U11199 ( .A(n31209), .B(net96340), .Y(n31220) );
  INVX1 U11200 ( .A(n31220), .Y(n23028) );
  AND2X1 U11201 ( .A(n31227), .B(net96340), .Y(n31234) );
  INVX1 U11202 ( .A(n31234), .Y(n23029) );
  AND2X2 U11203 ( .A(n29377), .B(n31229), .Y(n31240) );
  INVX1 U11204 ( .A(n31240), .Y(n23030) );
  INVX1 U11205 ( .A(n31240), .Y(n23031) );
  AND2X1 U11206 ( .A(n31249), .B(net96340), .Y(n31260) );
  INVX1 U11207 ( .A(n31260), .Y(n23032) );
  AND2X2 U11208 ( .A(n29378), .B(n31269), .Y(n31280) );
  INVX1 U11209 ( .A(n31280), .Y(n23034) );
  AND2X1 U11210 ( .A(n31287), .B(net96340), .Y(n31297) );
  AND2X1 U11211 ( .A(n31306), .B(net96340), .Y(n31316) );
  INVX1 U11212 ( .A(n31316), .Y(n23035) );
  AND2X1 U11213 ( .A(n31343), .B(net96340), .Y(n31354) );
  INVX1 U11214 ( .A(n31354), .Y(n23037) );
  AND2X1 U11215 ( .A(n31363), .B(net96340), .Y(n31374) );
  INVX1 U11216 ( .A(n31374), .Y(n23038) );
  AND2X1 U11217 ( .A(n31383), .B(net96340), .Y(n31394) );
  INVX1 U11218 ( .A(n31394), .Y(n23039) );
  AND2X1 U11219 ( .A(n31403), .B(net96340), .Y(n31414) );
  INVX1 U11220 ( .A(n31414), .Y(n23040) );
  AND2X1 U11221 ( .A(n31424), .B(net96340), .Y(n31435) );
  INVX1 U11222 ( .A(n31435), .Y(n23041) );
  INVX1 U11223 ( .A(n31454), .Y(n23042) );
  AND2X1 U11224 ( .A(n31463), .B(net96340), .Y(n31474) );
  INVX1 U11225 ( .A(n31474), .Y(n23043) );
  AND2X1 U11226 ( .A(n31483), .B(net96340), .Y(n31493) );
  AND2X1 U11227 ( .A(n31520), .B(net96340), .Y(n31531) );
  INVX1 U11228 ( .A(n31531), .Y(n23044) );
  AND2X1 U11229 ( .A(n31540), .B(net96340), .Y(n31551) );
  INVX1 U11230 ( .A(n31551), .Y(n23045) );
  AND2X1 U11231 ( .A(n31581), .B(net96340), .Y(n31592) );
  AND2X1 U11232 ( .A(n31601), .B(net96340), .Y(n31611) );
  INVX1 U11233 ( .A(n31611), .Y(n23046) );
  AND2X2 U11234 ( .A(n29374), .B(n31620), .Y(n31630) );
  INVX1 U11235 ( .A(n31630), .Y(n23047) );
  INVX1 U11236 ( .A(n31630), .Y(n23048) );
  AND2X1 U11237 ( .A(n31638), .B(net96340), .Y(n31647) );
  INVX1 U11238 ( .A(n31647), .Y(n23049) );
  AND2X2 U11239 ( .A(n20958), .B(n31656), .Y(n31667) );
  INVX1 U11240 ( .A(n31667), .Y(n23051) );
  INVX1 U11241 ( .A(n31667), .Y(n23052) );
  INVX1 U11242 ( .A(n31686), .Y(n23053) );
  AND2X1 U11243 ( .A(n31692), .B(net96340), .Y(n31699) );
  INVX1 U11244 ( .A(n31699), .Y(n23054) );
  AND2X2 U11245 ( .A(n29376), .B(n31694), .Y(n31705) );
  INVX1 U11246 ( .A(n31705), .Y(n23055) );
  INVX1 U11247 ( .A(n31705), .Y(n23056) );
  AND2X2 U11248 ( .A(n29376), .B(n31734), .Y(n31744) );
  INVX1 U11249 ( .A(n31744), .Y(n23057) );
  INVX1 U11250 ( .A(n31744), .Y(n23058) );
  AND2X1 U11251 ( .A(n31752), .B(net96340), .Y(n31763) );
  INVX1 U11252 ( .A(n31763), .Y(n23059) );
  AND2X2 U11253 ( .A(n29377), .B(n31772), .Y(n31783) );
  INVX1 U11254 ( .A(n31783), .Y(n23060) );
  AND2X1 U11255 ( .A(n31809), .B(net96340), .Y(n31816) );
  INVX1 U11256 ( .A(n31816), .Y(n23062) );
  AND2X2 U11257 ( .A(n31811), .B(n29375), .Y(n31822) );
  INVX1 U11258 ( .A(n31822), .Y(n23063) );
  INVX1 U11259 ( .A(n31822), .Y(n23064) );
  AND2X1 U11260 ( .A(n31831), .B(net96340), .Y(n31842) );
  INVX1 U11261 ( .A(n31842), .Y(n23065) );
  AND2X2 U11262 ( .A(n20957), .B(n31850), .Y(n31861) );
  INVX1 U11263 ( .A(n31861), .Y(n23066) );
  AND2X2 U11264 ( .A(n31871), .B(net96340), .Y(n31883) );
  AND2X2 U11265 ( .A(locTrig[1]), .B(n23206), .Y(n30635) );
  INVX1 U11266 ( .A(n30635), .Y(n23067) );
  AND2X2 U11267 ( .A(T[1]), .B(n21559), .Y(n33089) );
  INVX1 U11268 ( .A(n33089), .Y(n23068) );
  INVX1 U11269 ( .A(n33089), .Y(n23069) );
  AND2X2 U11270 ( .A(n25725), .B(n25327), .Y(n34266) );
  INVX1 U11271 ( .A(n34266), .Y(n23070) );
  INVX1 U11272 ( .A(n34266), .Y(n23071) );
  AND2X2 U11273 ( .A(n34302), .B(n25325), .Y(n34325) );
  INVX1 U11274 ( .A(n34325), .Y(n23072) );
  INVX1 U11275 ( .A(n34325), .Y(n23073) );
  AND2X2 U11276 ( .A(n25727), .B(pLoc[1]), .Y(n26061) );
  INVX1 U11277 ( .A(n26061), .Y(n23074) );
  INVX1 U11278 ( .A(n26061), .Y(n23075) );
  AND2X2 U11279 ( .A(n29376), .B(n30641), .Y(n30658) );
  INVX1 U11280 ( .A(n30658), .Y(n23076) );
  AND2X2 U11281 ( .A(n29381), .B(n30875), .Y(n30888) );
  INVX1 U11282 ( .A(n30888), .Y(n23077) );
  INVX1 U11283 ( .A(n30888), .Y(n23078) );
  AND2X2 U11284 ( .A(n20957), .B(n30977), .Y(n30989) );
  INVX1 U11285 ( .A(n30989), .Y(n23079) );
  AND2X2 U11286 ( .A(n34441), .B(n25714), .Y(n34349) );
  AND2X2 U11287 ( .A(direction_line[2]), .B(net145295), .Y(net95480) );
  INVX1 U11288 ( .A(net95480), .Y(net142788) );
  INVX1 U11289 ( .A(net95480), .Y(net142789) );
  BUFX2 U11290 ( .A(n25528), .Y(n23080) );
  AND2X2 U11291 ( .A(n25466), .B(n31286), .Y(n31298) );
  INVX1 U11292 ( .A(n31298), .Y(n23081) );
  INVX1 U11293 ( .A(n31298), .Y(n23082) );
  INVX1 U11294 ( .A(n25515), .Y(n23083) );
  INVX1 U11295 ( .A(n25515), .Y(n23084) );
  AND2X2 U11296 ( .A(n21527), .B(n29577), .Y(n13707) );
  INVX1 U11297 ( .A(n13707), .Y(n23085) );
  BUFX2 U11298 ( .A(n33064), .Y(n23086) );
  AND2X1 U11299 ( .A(n31893), .B(net96340), .Y(n24988) );
  INVX1 U11300 ( .A(n24988), .Y(n23087) );
  INVX1 U11301 ( .A(n21159), .Y(n23088) );
  BUFX2 U11302 ( .A(n33081), .Y(n26072) );
  AND2X2 U11303 ( .A(n34387), .B(n22988), .Y(n25653) );
  AND2X2 U11304 ( .A(n29377), .B(n31169), .Y(n31181) );
  INVX1 U11305 ( .A(n31181), .Y(n23089) );
  INVX1 U11306 ( .A(n31181), .Y(n23090) );
  BUFX2 U11307 ( .A(n15186), .Y(n23091) );
  AND2X2 U11308 ( .A(n29902), .B(n21106), .Y(n29803) );
  INVX1 U11309 ( .A(n29803), .Y(n23092) );
  AND2X2 U11310 ( .A(T[0]), .B(n33062), .Y(n33111) );
  AND2X2 U11311 ( .A(n33061), .B(n25679), .Y(n33066) );
  INVX1 U11312 ( .A(n33066), .Y(n23094) );
  INVX1 U11313 ( .A(n33066), .Y(n23095) );
  AND2X2 U11314 ( .A(n25336), .B(n22991), .Y(n33115) );
  INVX1 U11315 ( .A(n33115), .Y(n23096) );
  INVX1 U11316 ( .A(n33115), .Y(n23097) );
  AND2X2 U11317 ( .A(n33146), .B(n33105), .Y(n33107) );
  INVX1 U11318 ( .A(n33107), .Y(n23098) );
  INVX1 U11319 ( .A(n33107), .Y(n23099) );
  AND2X2 U11320 ( .A(n23296), .B(n29330), .Y(n32489) );
  INVX1 U11321 ( .A(n32489), .Y(n23100) );
  INVX1 U11322 ( .A(n32489), .Y(n23101) );
  AND2X2 U11323 ( .A(n29685), .B(n34503), .Y(n29584) );
  INVX1 U11324 ( .A(n29584), .Y(n23102) );
  INVX1 U11325 ( .A(n29584), .Y(n23103) );
  BUFX2 U11326 ( .A(n33143), .Y(n23104) );
  BUFX2 U11327 ( .A(n34253), .Y(n23105) );
  AND2X2 U11328 ( .A(n25688), .B(n25865), .Y(n25729) );
  AND2X2 U11329 ( .A(n2254), .B(n26050), .Y(n29475) );
  AND2X2 U11330 ( .A(n29510), .B(n26050), .Y(n29480) );
  INVX1 U11331 ( .A(n29480), .Y(n23106) );
  AND2X2 U11332 ( .A(n21236), .B(n21171), .Y(n34234) );
  BUFX2 U11333 ( .A(n29714), .Y(n23107) );
  BUFX2 U11334 ( .A(n29722), .Y(n23108) );
  BUFX2 U11335 ( .A(n29948), .Y(n23109) );
  AND2X2 U11336 ( .A(n23286), .B(n21106), .Y(n29760) );
  AND2X2 U11337 ( .A(n29835), .B(n30024), .Y(n33747) );
  AND2X2 U11338 ( .A(n30002), .B(n21106), .Y(n33560) );
  AND2X2 U11339 ( .A(n23298), .B(n32491), .Y(n32518) );
  OR2X2 U11340 ( .A(n22138), .B(n22110), .Y(n29846) );
  INVX1 U11341 ( .A(n29846), .Y(n23113) );
  INVX1 U11342 ( .A(n29846), .Y(n23114) );
  AND2X2 U11343 ( .A(n25466), .B(n31501), .Y(n31513) );
  INVX1 U11344 ( .A(n31513), .Y(n23115) );
  INVX1 U11345 ( .A(n31512), .Y(n23116) );
  AND2X2 U11346 ( .A(n23209), .B(n30795), .Y(n30808) );
  INVX1 U11347 ( .A(n30808), .Y(n23117) );
  INVX1 U11348 ( .A(n30808), .Y(n23118) );
  AND2X2 U11349 ( .A(n20966), .B(n30916), .Y(n30929) );
  INVX1 U11350 ( .A(n30929), .Y(n23119) );
  AND2X2 U11351 ( .A(n29378), .B(n30956), .Y(n30969) );
  INVX1 U11352 ( .A(n30969), .Y(n23120) );
  INVX1 U11353 ( .A(n30969), .Y(n23121) );
  AND2X2 U11354 ( .A(n20958), .B(n31131), .Y(n31144) );
  INVX1 U11355 ( .A(n31144), .Y(n23122) );
  AND2X2 U11356 ( .A(n25466), .B(n31342), .Y(n31355) );
  INVX1 U11357 ( .A(n31355), .Y(n23123) );
  INVX1 U11358 ( .A(n31355), .Y(n23124) );
  AND2X2 U11359 ( .A(n29378), .B(n31362), .Y(n31375) );
  INVX1 U11360 ( .A(n31375), .Y(n23125) );
  INVX1 U11361 ( .A(n31375), .Y(n23126) );
  AND2X2 U11362 ( .A(n29377), .B(n31580), .Y(n31593) );
  INVX1 U11363 ( .A(n31593), .Y(n23127) );
  INVX1 U11364 ( .A(n31593), .Y(n23128) );
  AND2X2 U11365 ( .A(n25466), .B(n31791), .Y(n31804) );
  INVX1 U11366 ( .A(n31804), .Y(n23129) );
  INVX1 U11367 ( .A(n31804), .Y(n23130) );
  AND2X2 U11368 ( .A(n29378), .B(n31830), .Y(n31843) );
  INVX1 U11369 ( .A(n31843), .Y(n23131) );
  INVX1 U11370 ( .A(n31843), .Y(n23132) );
  AND2X2 U11371 ( .A(n27074), .B(n25644), .Y(n34312) );
  AND2X2 U11372 ( .A(n25833), .B(n25201), .Y(n34433) );
  AND2X2 U11373 ( .A(n29381), .B(n30895), .Y(n30908) );
  INVX1 U11374 ( .A(n30908), .Y(n23133) );
  INVX1 U11375 ( .A(n30908), .Y(n23134) );
  AND2X2 U11376 ( .A(n25466), .B(n31382), .Y(n31395) );
  INVX1 U11377 ( .A(n31395), .Y(n23135) );
  INVX1 U11378 ( .A(n31395), .Y(n23136) );
  AND2X2 U11379 ( .A(n29377), .B(n31462), .Y(n31475) );
  INVX1 U11380 ( .A(n31475), .Y(n23137) );
  INVX1 U11381 ( .A(n31475), .Y(n23138) );
  BUFX2 U11382 ( .A(n33109), .Y(n23139) );
  OR2X2 U11383 ( .A(n8037), .B(n8036), .Y(n29502) );
  INVX1 U11384 ( .A(n29502), .Y(n23140) );
  AND2X2 U11385 ( .A(net146838), .B(net143010), .Y(n25130) );
  INVX1 U11386 ( .A(n25130), .Y(n23141) );
  INVX1 U11387 ( .A(n25130), .Y(n23142) );
  AND2X2 U11388 ( .A(n29565), .B(n29564), .Y(n29570) );
  INVX1 U11389 ( .A(n29570), .Y(n23143) );
  INVX1 U11390 ( .A(n29570), .Y(n23144) );
  AND2X2 U11391 ( .A(n29376), .B(n30672), .Y(n30688) );
  INVX1 U11392 ( .A(n30688), .Y(n23145) );
  INVX1 U11393 ( .A(n30688), .Y(n23146) );
  AND2X2 U11394 ( .A(n29378), .B(n30695), .Y(n30708) );
  INVX1 U11395 ( .A(n30708), .Y(n23147) );
  INVX1 U11396 ( .A(n30708), .Y(n23148) );
  AND2X2 U11397 ( .A(n29381), .B(n30715), .Y(n30728) );
  INVX1 U11398 ( .A(n30728), .Y(n23149) );
  AND2X2 U11399 ( .A(n29381), .B(n30734), .Y(n30747) );
  INVX1 U11400 ( .A(n30747), .Y(n23150) );
  AND2X2 U11401 ( .A(n29381), .B(n30755), .Y(n30768) );
  INVX1 U11402 ( .A(n30768), .Y(n23151) );
  INVX1 U11403 ( .A(n30768), .Y(n23152) );
  AND2X2 U11404 ( .A(n29381), .B(n30774), .Y(n30787) );
  INVX1 U11405 ( .A(n30787), .Y(n23153) );
  INVX1 U11406 ( .A(n30787), .Y(n23154) );
  AND2X2 U11407 ( .A(n29381), .B(n30814), .Y(n30827) );
  INVX1 U11408 ( .A(n30827), .Y(n23155) );
  INVX1 U11409 ( .A(n30827), .Y(n23156) );
  AND2X2 U11410 ( .A(n29381), .B(n30854), .Y(n30867) );
  INVX1 U11411 ( .A(n30867), .Y(n23157) );
  AND2X2 U11412 ( .A(n29376), .B(n31013), .Y(n31026) );
  INVX1 U11413 ( .A(n31026), .Y(n23158) );
  INVX1 U11414 ( .A(n31026), .Y(n23159) );
  AND2X2 U11415 ( .A(n20966), .B(n31051), .Y(n31064) );
  INVX1 U11416 ( .A(n31064), .Y(n23160) );
  INVX1 U11417 ( .A(n31064), .Y(n23161) );
  AND2X2 U11418 ( .A(n29376), .B(n31091), .Y(n31104) );
  INVX1 U11419 ( .A(n31104), .Y(n23162) );
  INVX1 U11420 ( .A(n31104), .Y(n23163) );
  AND2X2 U11421 ( .A(n23209), .B(n31208), .Y(n31221) );
  INVX1 U11422 ( .A(n31221), .Y(n23164) );
  INVX1 U11423 ( .A(n31221), .Y(n23165) );
  AND2X2 U11424 ( .A(n25466), .B(n31248), .Y(n31261) );
  INVX1 U11425 ( .A(n31261), .Y(n23166) );
  INVX1 U11426 ( .A(n31261), .Y(n23167) );
  AND2X2 U11427 ( .A(n29376), .B(n31402), .Y(n31415) );
  INVX1 U11428 ( .A(n31415), .Y(n23168) );
  INVX1 U11429 ( .A(n31415), .Y(n23169) );
  AND2X2 U11430 ( .A(n25466), .B(n31423), .Y(n31436) );
  INVX1 U11431 ( .A(n31436), .Y(n23170) );
  INVX1 U11432 ( .A(n31436), .Y(n23171) );
  AND2X2 U11433 ( .A(n25466), .B(n31443), .Y(n31455) );
  INVX1 U11434 ( .A(n31455), .Y(n23172) );
  INVX1 U11435 ( .A(n31455), .Y(n23173) );
  AND2X2 U11436 ( .A(n29378), .B(n31519), .Y(n31532) );
  INVX1 U11437 ( .A(n31532), .Y(n23174) );
  INVX1 U11438 ( .A(n31532), .Y(n23175) );
  AND2X2 U11439 ( .A(n29377), .B(n31539), .Y(n31552) );
  INVX1 U11440 ( .A(n31552), .Y(n23176) );
  INVX1 U11441 ( .A(n31552), .Y(n23177) );
  AND2X2 U11442 ( .A(n29378), .B(n31559), .Y(n31572) );
  INVX1 U11443 ( .A(n31572), .Y(n23178) );
  INVX1 U11444 ( .A(n31572), .Y(n23179) );
  AND2X2 U11445 ( .A(n25466), .B(n31674), .Y(n31687) );
  INVX1 U11446 ( .A(n31687), .Y(n23180) );
  AND2X2 U11447 ( .A(n29376), .B(n31713), .Y(n31726) );
  INVX1 U11448 ( .A(n31726), .Y(n23181) );
  INVX1 U11449 ( .A(n31726), .Y(n23182) );
  AND2X2 U11450 ( .A(n29377), .B(n31751), .Y(n31764) );
  INVX1 U11451 ( .A(n31764), .Y(n23183) );
  INVX1 U11452 ( .A(n31764), .Y(n23184) );
  AND2X2 U11453 ( .A(n29376), .B(n31870), .Y(n31884) );
  INVX1 U11454 ( .A(n31884), .Y(n23185) );
  INVX1 U11455 ( .A(n31884), .Y(n23186) );
  AND2X2 U11456 ( .A(n34237), .B(n23000), .Y(n34252) );
  INVX1 U11457 ( .A(n34252), .Y(n23187) );
  BUFX2 U11458 ( .A(n33137), .Y(n23188) );
  INVX1 U11459 ( .A(n30687), .Y(n23189) );
  AND2X2 U11460 ( .A(n29381), .B(n30835), .Y(n30848) );
  INVX1 U11461 ( .A(n30848), .Y(n23190) );
  INVX1 U11462 ( .A(n30848), .Y(n23191) );
  INVX1 U11463 ( .A(n30866), .Y(n23192) );
  AND2X2 U11464 ( .A(n29372), .B(n21553), .Y(n30948) );
  INVX1 U11465 ( .A(n30948), .Y(n23193) );
  INVX1 U11466 ( .A(n30948), .Y(n23194) );
  INVX1 U11467 ( .A(n31025), .Y(n23195) );
  INVX1 U11468 ( .A(n31103), .Y(n23196) );
  AND2X2 U11469 ( .A(n29376), .B(n31322), .Y(n31335) );
  INVX1 U11470 ( .A(n31335), .Y(n23197) );
  INVX1 U11471 ( .A(n31335), .Y(n23198) );
  INVX1 U11472 ( .A(n31571), .Y(n23199) );
  BUFX2 U11473 ( .A(n30651), .Y(n23200) );
  BUFX2 U11474 ( .A(net95464), .Y(net142478) );
  BUFX2 U11475 ( .A(n25648), .Y(n23201) );
  BUFX2 U11476 ( .A(n25640), .Y(n23202) );
  AND2X2 U11477 ( .A(n25485), .B(n25621), .Y(n25859) );
  BUFX2 U11478 ( .A(n34316), .Y(n23203) );
  BUFX2 U11479 ( .A(n29727), .Y(n23204) );
  BUFX2 U11480 ( .A(grid[331]), .Y(n23205) );
  AND2X2 U11481 ( .A(n29484), .B(n25589), .Y(n23206) );
  MUX2X1 U11482 ( .B(n25516), .A(grid[97]), .S(n21091), .Y(n28324) );
  INVX2 U11483 ( .A(n26514), .Y(n26504) );
  OR2X2 U11484 ( .A(net109469), .B(n4225), .Y(n23207) );
  INVX1 U11485 ( .A(n30045), .Y(n29503) );
  INVX1 U11486 ( .A(n26446), .Y(n23208) );
  INVX1 U11487 ( .A(n30675), .Y(n23212) );
  INVX1 U11488 ( .A(n30677), .Y(n23213) );
  INVX1 U11489 ( .A(n30698), .Y(n23215) );
  INVX1 U11490 ( .A(n30700), .Y(n23216) );
  INVX1 U11491 ( .A(n30718), .Y(n23218) );
  INVX1 U11492 ( .A(n30720), .Y(n23219) );
  INVX1 U11493 ( .A(n30737), .Y(n23221) );
  INVX1 U11494 ( .A(n30739), .Y(n23222) );
  INVX1 U11495 ( .A(n30758), .Y(n23224) );
  INVX1 U11496 ( .A(n30760), .Y(n23225) );
  INVX1 U11497 ( .A(n30777), .Y(n23228) );
  INVX1 U11498 ( .A(n30779), .Y(n23229) );
  INVX1 U11499 ( .A(n30798), .Y(n23231) );
  INVX1 U11500 ( .A(n30800), .Y(n23232) );
  INVX1 U11501 ( .A(n30817), .Y(n23235) );
  INVX1 U11502 ( .A(n30819), .Y(n23236) );
  INVX1 U11503 ( .A(n30857), .Y(n23238) );
  INVX1 U11504 ( .A(n30859), .Y(n23239) );
  INVX1 U11505 ( .A(n30919), .Y(n23241) );
  INVX1 U11506 ( .A(n30921), .Y(n23242) );
  INVX1 U11507 ( .A(n31094), .Y(n23244) );
  INVX1 U11508 ( .A(n31096), .Y(n23245) );
  INVX1 U11509 ( .A(n31211), .Y(n23247) );
  INVX1 U11510 ( .A(n31213), .Y(n23248) );
  INVX1 U11511 ( .A(n31251), .Y(n23250) );
  INVX1 U11512 ( .A(n31253), .Y(n23251) );
  INVX1 U11513 ( .A(n31503), .Y(n23253) );
  INVX1 U11514 ( .A(n31505), .Y(n23254) );
  INVX1 U11515 ( .A(n31542), .Y(n23256) );
  INVX1 U11516 ( .A(n31544), .Y(n23257) );
  INVX1 U11517 ( .A(n31562), .Y(n23260) );
  INVX1 U11518 ( .A(n31564), .Y(n23261) );
  INVX1 U11519 ( .A(n31677), .Y(n23263) );
  INVX1 U11520 ( .A(n31679), .Y(n23264) );
  INVX1 U11521 ( .A(n31716), .Y(n23267) );
  INVX1 U11522 ( .A(n31718), .Y(n23268) );
  INVX1 U11523 ( .A(n31910), .Y(n23270) );
  INVX1 U11524 ( .A(n21042), .Y(n23271) );
  AND2X2 U11525 ( .A(n25426), .B(n25452), .Y(n23273) );
  AND2X2 U11526 ( .A(n33056), .B(n33055), .Y(n23274) );
  AND2X2 U11527 ( .A(n29835), .B(n29943), .Y(n23275) );
  AND2X2 U11528 ( .A(n29352), .B(net96340), .Y(n23276) );
  OR2X2 U11529 ( .A(n25681), .B(n25320), .Y(n23277) );
  OR2X2 U11530 ( .A(net109417), .B(net150331), .Y(net138174) );
  AND2X2 U11531 ( .A(n29725), .B(n29726), .Y(n23278) );
  AND2X2 U11532 ( .A(net110927), .B(net150330), .Y(n23279) );
  AND2X2 U11533 ( .A(states[1]), .B(n20972), .Y(n23280) );
  AND2X2 U11534 ( .A(wT), .B(n27117), .Y(n23281) );
  AND2X2 U11535 ( .A(n29724), .B(n29191), .Y(net138161) );
  AND2X2 U11536 ( .A(n29811), .B(n27313), .Y(n23282) );
  AND2X2 U11537 ( .A(n30012), .B(n27313), .Y(n23283) );
  AND2X2 U11538 ( .A(n29925), .B(n27314), .Y(n23284) );
  AND2X2 U11539 ( .A(n27294), .B(n29825), .Y(n23285) );
  AND2X2 U11540 ( .A(n27313), .B(n29831), .Y(n23286) );
  AND2X2 U11541 ( .A(n27103), .B(n25332), .Y(n23287) );
  AND2X2 U11542 ( .A(n27294), .B(n29811), .Y(n23288) );
  AND2X2 U11543 ( .A(n27313), .B(n29815), .Y(n23289) );
  AND2X2 U11544 ( .A(n27294), .B(n30012), .Y(n23290) );
  AND2X2 U11545 ( .A(n27313), .B(n29925), .Y(n23291) );
  AND2X2 U11546 ( .A(n27021), .B(n32773), .Y(n23292) );
  AND2X2 U11547 ( .A(n27294), .B(n29831), .Y(n23293) );
  AND2X2 U11548 ( .A(n27313), .B(n29967), .Y(n23294) );
  AND2X2 U11549 ( .A(n27294), .B(n29815), .Y(n23295) );
  AND2X2 U11550 ( .A(n27314), .B(n21211), .Y(n23296) );
  AND2X2 U11551 ( .A(n30012), .B(n27315), .Y(n23297) );
  AND2X2 U11552 ( .A(n27294), .B(n29925), .Y(n23298) );
  AND2X2 U11553 ( .A(n27313), .B(n21211), .Y(n23299) );
  AND2X2 U11554 ( .A(n26942), .B(n25147), .Y(n23300) );
  AND2X2 U11555 ( .A(n29825), .B(n27313), .Y(n23301) );
  AND2X2 U11556 ( .A(n33682), .B(n25148), .Y(n23302) );
  AND2X2 U11557 ( .A(n27207), .B(n25149), .Y(n23303) );
  AND2X2 U11558 ( .A(n25424), .B(n26078), .Y(n23304) );
  AND2X2 U11559 ( .A(n25403), .B(n25202), .Y(n23305) );
  AND2X2 U11560 ( .A(n29922), .B(n29330), .Y(n23306) );
  AND2X2 U11561 ( .A(n29933), .B(n29330), .Y(n23307) );
  AND2X2 U11562 ( .A(n26879), .B(n27195), .Y(n23308) );
  AND2X2 U11563 ( .A(n24979), .B(n22989), .Y(n23309) );
  AND2X2 U11564 ( .A(n27265), .B(n27239), .Y(n23310) );
  AND2X2 U11565 ( .A(n27238), .B(n27222), .Y(n23311) );
  AND2X2 U11566 ( .A(n27238), .B(n27240), .Y(n23312) );
  AND2X2 U11567 ( .A(n27238), .B(n30434), .Y(n23313) );
  AND2X2 U11568 ( .A(n27238), .B(n30443), .Y(n23314) );
  AND2X2 U11569 ( .A(n27238), .B(n30451), .Y(n23315) );
  AND2X2 U11570 ( .A(n27238), .B(n23613), .Y(n23316) );
  AND2X2 U11571 ( .A(n27238), .B(n30465), .Y(n23317) );
  AND2X2 U11572 ( .A(n27270), .B(n27222), .Y(n23318) );
  AND2X2 U11573 ( .A(n27270), .B(n27240), .Y(n23319) );
  AND2X2 U11574 ( .A(n27270), .B(n30434), .Y(n23320) );
  AND2X2 U11575 ( .A(n27306), .B(n23442), .Y(n23321) );
  AND2X2 U11576 ( .A(n27270), .B(n30443), .Y(n23322) );
  AND2X2 U11577 ( .A(n27270), .B(n30451), .Y(n23323) );
  AND2X2 U11578 ( .A(n27270), .B(n23613), .Y(n23324) );
  AND2X2 U11579 ( .A(n27270), .B(n30473), .Y(n23325) );
  AND2X2 U11580 ( .A(n30226), .B(n26163), .Y(n23326) );
  AND2X2 U11581 ( .A(n30227), .B(n27239), .Y(n23327) );
  AND2X2 U11582 ( .A(n30228), .B(n27222), .Y(n23328) );
  AND2X2 U11583 ( .A(n30226), .B(n27268), .Y(n23329) );
  AND2X2 U11584 ( .A(n30228), .B(n27240), .Y(n23330) );
  AND2X2 U11585 ( .A(n30226), .B(n21405), .Y(n23331) );
  AND2X2 U11586 ( .A(n30227), .B(n30433), .Y(n23332) );
  AND2X2 U11587 ( .A(n30228), .B(n30434), .Y(n23333) );
  AND2X2 U11588 ( .A(n30226), .B(n23442), .Y(n23334) );
  AND2X2 U11589 ( .A(n30228), .B(n30443), .Y(n23335) );
  AND2X2 U11590 ( .A(n30227), .B(n30450), .Y(n23336) );
  AND2X2 U11591 ( .A(n30228), .B(n30451), .Y(n23337) );
  AND2X2 U11592 ( .A(n30226), .B(n27308), .Y(n23338) );
  AND2X2 U11593 ( .A(n30228), .B(n23613), .Y(n23339) );
  AND2X2 U11594 ( .A(n30227), .B(n30464), .Y(n23340) );
  AND2X2 U11595 ( .A(n30228), .B(n30465), .Y(n23341) );
  AND2X2 U11596 ( .A(n30226), .B(n30410), .Y(n23342) );
  AND2X2 U11597 ( .A(n30228), .B(n30473), .Y(n23343) );
  AND2X2 U11598 ( .A(n30273), .B(n27239), .Y(n23344) );
  AND2X2 U11599 ( .A(n30274), .B(n27222), .Y(n23345) );
  AND2X2 U11600 ( .A(n21414), .B(n27268), .Y(n23346) );
  AND2X2 U11601 ( .A(n30273), .B(n30433), .Y(n23347) );
  AND2X2 U11602 ( .A(n30274), .B(n30434), .Y(n23348) );
  AND2X2 U11603 ( .A(n21414), .B(n23442), .Y(n23349) );
  AND2X2 U11604 ( .A(n30274), .B(n30443), .Y(n23350) );
  AND2X2 U11605 ( .A(n30273), .B(n30450), .Y(n23351) );
  AND2X2 U11606 ( .A(n30274), .B(n30451), .Y(n23352) );
  AND2X2 U11607 ( .A(n21414), .B(n27308), .Y(n23353) );
  AND2X2 U11608 ( .A(n30274), .B(n23613), .Y(n23354) );
  AND2X2 U11609 ( .A(n30273), .B(n30464), .Y(n23355) );
  AND2X2 U11610 ( .A(n30274), .B(n30465), .Y(n23356) );
  AND2X2 U11611 ( .A(n30274), .B(n30473), .Y(n23357) );
  AND2X2 U11612 ( .A(n30320), .B(n27239), .Y(n23358) );
  AND2X2 U11613 ( .A(n30321), .B(n27222), .Y(n23359) );
  AND2X2 U11614 ( .A(n30320), .B(n27237), .Y(n23360) );
  AND2X2 U11615 ( .A(n30321), .B(n27240), .Y(n23361) );
  AND2X2 U11616 ( .A(n30320), .B(n30433), .Y(n23362) );
  AND2X2 U11617 ( .A(n30321), .B(n30434), .Y(n23363) );
  AND2X2 U11618 ( .A(n27266), .B(n23442), .Y(n23364) );
  AND2X2 U11619 ( .A(n30320), .B(n30442), .Y(n23365) );
  AND2X2 U11620 ( .A(n30321), .B(n30443), .Y(n23366) );
  AND2X2 U11621 ( .A(n30320), .B(n30450), .Y(n23367) );
  AND2X2 U11622 ( .A(n30321), .B(n30451), .Y(n23368) );
  AND2X2 U11623 ( .A(n30320), .B(n30458), .Y(n23369) );
  AND2X2 U11624 ( .A(n30321), .B(n23613), .Y(n23370) );
  AND2X2 U11625 ( .A(n30320), .B(n30464), .Y(n23371) );
  AND2X2 U11626 ( .A(n30321), .B(n30465), .Y(n23372) );
  AND2X2 U11627 ( .A(n30320), .B(n30476), .Y(n23373) );
  AND2X2 U11628 ( .A(n30321), .B(n30473), .Y(n23374) );
  AND2X2 U11629 ( .A(n30364), .B(n27239), .Y(n23375) );
  AND2X2 U11630 ( .A(n30365), .B(n27222), .Y(n23376) );
  AND2X2 U11631 ( .A(n30364), .B(n27237), .Y(n23377) );
  AND2X2 U11632 ( .A(n30365), .B(n27240), .Y(n23378) );
  AND2X2 U11633 ( .A(n30364), .B(n30433), .Y(n23379) );
  AND2X2 U11634 ( .A(n30365), .B(n30434), .Y(n23380) );
  AND2X2 U11635 ( .A(n27305), .B(n23442), .Y(n23381) );
  AND2X2 U11636 ( .A(n30364), .B(n30442), .Y(n23382) );
  AND2X2 U11637 ( .A(n30365), .B(n30443), .Y(n23383) );
  AND2X2 U11638 ( .A(n30364), .B(n30450), .Y(n23384) );
  AND2X2 U11639 ( .A(n30365), .B(n30451), .Y(n23385) );
  AND2X2 U11640 ( .A(n30364), .B(n30458), .Y(n23386) );
  AND2X2 U11641 ( .A(n30365), .B(n23613), .Y(n23387) );
  AND2X2 U11642 ( .A(n30364), .B(n30464), .Y(n23388) );
  AND2X2 U11643 ( .A(n30365), .B(n30465), .Y(n23389) );
  AND2X2 U11644 ( .A(n30364), .B(n30476), .Y(n23390) );
  AND2X2 U11645 ( .A(n30365), .B(n30473), .Y(n23391) );
  AND2X2 U11646 ( .A(n30411), .B(n27239), .Y(n23392) );
  AND2X2 U11647 ( .A(n30412), .B(n27222), .Y(n23393) );
  AND2X2 U11648 ( .A(n27264), .B(n27268), .Y(n23394) );
  AND2X2 U11649 ( .A(n30412), .B(n27240), .Y(n23395) );
  AND2X2 U11650 ( .A(n30411), .B(n30433), .Y(n23396) );
  AND2X2 U11651 ( .A(n30412), .B(n30434), .Y(n23397) );
  AND2X2 U11652 ( .A(n27264), .B(n23442), .Y(n23398) );
  AND2X2 U11653 ( .A(n30412), .B(n30443), .Y(n23399) );
  AND2X2 U11654 ( .A(n30411), .B(n30450), .Y(n23400) );
  AND2X2 U11655 ( .A(n30412), .B(n30451), .Y(n23401) );
  AND2X2 U11656 ( .A(n27264), .B(n27308), .Y(n23402) );
  AND2X2 U11657 ( .A(n30412), .B(n23613), .Y(n23403) );
  AND2X2 U11658 ( .A(n30411), .B(n30464), .Y(n23404) );
  AND2X2 U11659 ( .A(n30412), .B(n30465), .Y(n23405) );
  AND2X2 U11660 ( .A(n27264), .B(n30410), .Y(n23406) );
  AND2X2 U11661 ( .A(n30476), .B(n30411), .Y(n23407) );
  AND2X2 U11662 ( .A(n30473), .B(n30412), .Y(n23408) );
  AND2X2 U11663 ( .A(n27239), .B(n30475), .Y(n23409) );
  AND2X2 U11664 ( .A(n27222), .B(n30472), .Y(n23410) );
  AND2X2 U11665 ( .A(n27268), .B(n29670), .Y(n23411) );
  AND2X2 U11666 ( .A(n27240), .B(n30472), .Y(n23412) );
  AND2X2 U11667 ( .A(n30433), .B(n30475), .Y(n23413) );
  AND2X2 U11668 ( .A(n30434), .B(n30472), .Y(n23414) );
  AND2X2 U11669 ( .A(n23442), .B(n29670), .Y(n23415) );
  AND2X2 U11670 ( .A(n30443), .B(n30472), .Y(n23416) );
  AND2X2 U11671 ( .A(n30450), .B(n30475), .Y(n23417) );
  AND2X2 U11672 ( .A(n30451), .B(n30472), .Y(n23418) );
  AND2X2 U11673 ( .A(n27308), .B(n29670), .Y(n23419) );
  AND2X2 U11674 ( .A(n30458), .B(n30475), .Y(n23420) );
  AND2X2 U11675 ( .A(n23613), .B(n30472), .Y(n23421) );
  AND2X2 U11676 ( .A(n30464), .B(n30475), .Y(n23422) );
  AND2X2 U11677 ( .A(n30465), .B(n30472), .Y(n23423) );
  AND2X2 U11678 ( .A(n27198), .B(n25115), .Y(n23424) );
  INVX2 U11679 ( .A(n32197), .Y(n29319) );
  AND2X2 U11680 ( .A(n34174), .B(n23443), .Y(n23425) );
  AND2X2 U11681 ( .A(n24324), .B(n25204), .Y(n23426) );
  AND2X2 U11682 ( .A(n25855), .B(n23093), .Y(n23427) );
  AND2X2 U11683 ( .A(n29191), .B(net96340), .Y(n23428) );
  INVX1 U11684 ( .A(n33262), .Y(n23429) );
  INVX1 U11685 ( .A(n23429), .Y(n23430) );
  INVX1 U11686 ( .A(n34359), .Y(n23431) );
  INVX1 U11687 ( .A(n23431), .Y(n23432) );
  INVX1 U11688 ( .A(n33007), .Y(n23433) );
  INVX1 U11689 ( .A(n23433), .Y(n23434) );
  AND2X2 U11690 ( .A(n3246), .B(n33326), .Y(n32542) );
  INVX1 U11691 ( .A(n32542), .Y(n23435) );
  INVX1 U11692 ( .A(n32543), .Y(n23436) );
  INVX1 U11693 ( .A(n23436), .Y(n23437) );
  AND2X2 U11694 ( .A(n22982), .B(n25842), .Y(n31484) );
  INVX1 U11695 ( .A(n31484), .Y(n23438) );
  AND2X2 U11696 ( .A(n23128), .B(n25182), .Y(n31582) );
  INVX1 U11697 ( .A(n31582), .Y(n23439) );
  BUFX2 U11698 ( .A(n29569), .Y(n34189) );
  INVX1 U11699 ( .A(n34189), .Y(n23440) );
  INVX1 U11700 ( .A(n34189), .Y(n23441) );
  INVX2 U11701 ( .A(n25110), .Y(n23442) );
  INVX1 U11702 ( .A(n29662), .Y(n30441) );
  AND2X2 U11703 ( .A(net90055), .B(n34338), .Y(n23443) );
  INVX1 U11704 ( .A(n25121), .Y(n23444) );
  INVX1 U11705 ( .A(n21372), .Y(n23445) );
  INVX1 U11706 ( .A(n21372), .Y(n23446) );
  INVX1 U11707 ( .A(n25124), .Y(n23447) );
  INVX1 U11708 ( .A(n21381), .Y(n23448) );
  INVX1 U11709 ( .A(n21381), .Y(n23449) );
  AND2X2 U11710 ( .A(n29943), .B(n21106), .Y(n23450) );
  AND2X2 U11711 ( .A(n23297), .B(n29331), .Y(n23451) );
  INVX1 U11712 ( .A(n21390), .Y(n23452) );
  INVX1 U11713 ( .A(n21390), .Y(n23453) );
  INVX1 U11714 ( .A(n21390), .Y(n23454) );
  INVX1 U11715 ( .A(n21390), .Y(n23455) );
  AND2X2 U11716 ( .A(n30274), .B(n27240), .Y(n23456) );
  AND2X2 U11717 ( .A(n30626), .B(n29922), .Y(n23457) );
  AND2X2 U11718 ( .A(n29225), .B(n26593), .Y(n30648) );
  INVX1 U11719 ( .A(n30648), .Y(n23458) );
  AND2X2 U11720 ( .A(n25882), .B(n32299), .Y(n31100) );
  INVX1 U11721 ( .A(n31100), .Y(n23459) );
  AND2X2 U11722 ( .A(n29223), .B(n26648), .Y(n31173) );
  INVX1 U11723 ( .A(n31173), .Y(n23460) );
  AND2X2 U11724 ( .A(n29223), .B(n26596), .Y(n31504) );
  AND2X2 U11725 ( .A(n29222), .B(n27163), .Y(n31523) );
  INVX1 U11726 ( .A(n31523), .Y(n23461) );
  AND2X2 U11727 ( .A(n29222), .B(n26862), .Y(n31603) );
  INVX1 U11728 ( .A(n31603), .Y(n23462) );
  AND2X2 U11729 ( .A(n29288), .B(n26975), .Y(n31628) );
  INVX1 U11730 ( .A(n31628), .Y(n23463) );
  INVX1 U11731 ( .A(n32589), .Y(n23464) );
  AND2X2 U11732 ( .A(n22987), .B(n23087), .Y(n31909) );
  INVX1 U11733 ( .A(net111600), .Y(net137830) );
  INVX1 U11734 ( .A(n23092), .Y(n23466) );
  INVX8 U11735 ( .A(n25148), .Y(n23468) );
  INVX8 U11736 ( .A(n25149), .Y(n23469) );
  AND2X2 U11737 ( .A(n23294), .B(n25723), .Y(n23470) );
  INVX1 U11738 ( .A(n23101), .Y(n23471) );
  INVX1 U11739 ( .A(n23100), .Y(n32973) );
  INVX1 U11740 ( .A(n31554), .Y(n23472) );
  MUX2X1 U11741 ( .B(n28507), .A(n28508), .S(n26491), .Y(n28506) );
  AND2X2 U11742 ( .A(n33045), .B(n33044), .Y(n33046) );
  AND2X2 U11743 ( .A(n3239), .B(n25680), .Y(n23473) );
  AND2X2 U11744 ( .A(n3233), .B(n25657), .Y(n23474) );
  AND2X2 U11745 ( .A(n29617), .B(n29616), .Y(n23475) );
  INVX1 U11746 ( .A(n33033), .Y(n25462) );
  INVX8 U11747 ( .A(n25661), .Y(n27911) );
  BUFX2 U11748 ( .A(n32971), .Y(n27175) );
  INVX1 U11749 ( .A(net112192), .Y(net137489) );
  INVX1 U11750 ( .A(n29499), .Y(n23476) );
  INVX1 U11751 ( .A(n23476), .Y(n23477) );
  BUFX2 U11752 ( .A(n29734), .Y(n23478) );
  BUFX2 U11753 ( .A(n29747), .Y(n23479) );
  BUFX2 U11754 ( .A(n30084), .Y(n23480) );
  BUFX2 U11755 ( .A(n30091), .Y(n23481) );
  BUFX2 U11756 ( .A(n30099), .Y(n23482) );
  BUFX2 U11757 ( .A(n30108), .Y(n23483) );
  BUFX2 U11758 ( .A(n30116), .Y(n23484) );
  BUFX2 U11759 ( .A(n30125), .Y(n23485) );
  BUFX2 U11760 ( .A(n30134), .Y(n23486) );
  BUFX2 U11761 ( .A(n30142), .Y(n23487) );
  BUFX2 U11762 ( .A(n30148), .Y(n23488) );
  BUFX2 U11763 ( .A(n30153), .Y(n23489) );
  BUFX2 U11764 ( .A(n30158), .Y(n23490) );
  BUFX2 U11765 ( .A(n30163), .Y(n23491) );
  BUFX2 U11766 ( .A(n30168), .Y(n23492) );
  BUFX2 U11767 ( .A(n30173), .Y(n23493) );
  BUFX2 U11768 ( .A(n30178), .Y(n23494) );
  BUFX2 U11769 ( .A(n30184), .Y(n23495) );
  BUFX2 U11770 ( .A(n30194), .Y(n23496) );
  BUFX2 U11771 ( .A(n30199), .Y(n23497) );
  BUFX2 U11772 ( .A(n30204), .Y(n23498) );
  BUFX2 U11773 ( .A(n30209), .Y(n23499) );
  BUFX2 U11774 ( .A(n30214), .Y(n23500) );
  BUFX2 U11775 ( .A(n30219), .Y(n23501) );
  BUFX2 U11776 ( .A(n30224), .Y(n23502) );
  BUFX2 U11777 ( .A(n30233), .Y(n23503) );
  BUFX2 U11778 ( .A(n30242), .Y(n23504) );
  BUFX2 U11779 ( .A(n30247), .Y(n23505) );
  BUFX2 U11780 ( .A(n30252), .Y(n23506) );
  BUFX2 U11781 ( .A(n30257), .Y(n23507) );
  BUFX2 U11782 ( .A(n30262), .Y(n23508) );
  BUFX2 U11783 ( .A(n30267), .Y(n23509) );
  BUFX2 U11784 ( .A(n30271), .Y(n23510) );
  BUFX2 U11785 ( .A(n30279), .Y(n23511) );
  BUFX2 U11786 ( .A(n30288), .Y(n23512) );
  BUFX2 U11787 ( .A(n30293), .Y(n23513) );
  BUFX2 U11788 ( .A(n30298), .Y(n23514) );
  BUFX2 U11789 ( .A(n30303), .Y(n23515) );
  BUFX2 U11790 ( .A(n30308), .Y(n23516) );
  BUFX2 U11791 ( .A(n30313), .Y(n23517) );
  BUFX2 U11792 ( .A(n30318), .Y(n23518) );
  BUFX2 U11793 ( .A(n30326), .Y(n23519) );
  BUFX2 U11794 ( .A(n30334), .Y(n23520) );
  BUFX2 U11795 ( .A(n30339), .Y(n23521) );
  BUFX2 U11796 ( .A(n30344), .Y(n23522) );
  BUFX2 U11797 ( .A(n30348), .Y(n23523) );
  BUFX2 U11798 ( .A(n30353), .Y(n23524) );
  BUFX2 U11799 ( .A(n30358), .Y(n23525) );
  BUFX2 U11800 ( .A(n30363), .Y(n23526) );
  BUFX2 U11801 ( .A(n30370), .Y(n23527) );
  BUFX2 U11802 ( .A(n30379), .Y(n23528) );
  BUFX2 U11803 ( .A(n30384), .Y(n23529) );
  BUFX2 U11804 ( .A(n30388), .Y(n23530) );
  BUFX2 U11805 ( .A(n30393), .Y(n23531) );
  BUFX2 U11806 ( .A(n30398), .Y(n23532) );
  BUFX2 U11807 ( .A(n30403), .Y(n23533) );
  BUFX2 U11808 ( .A(n30408), .Y(n23534) );
  BUFX2 U11809 ( .A(n30417), .Y(n23535) );
  BUFX2 U11810 ( .A(n30425), .Y(n23536) );
  BUFX2 U11811 ( .A(n30431), .Y(n23537) );
  BUFX2 U11812 ( .A(n30439), .Y(n23538) );
  BUFX2 U11813 ( .A(n30448), .Y(n23539) );
  BUFX2 U11814 ( .A(n30456), .Y(n23540) );
  BUFX2 U11815 ( .A(n30463), .Y(n23541) );
  BUFX2 U11816 ( .A(n30470), .Y(n23542) );
  BUFX2 U11817 ( .A(n33195), .Y(n23543) );
  INVX1 U11818 ( .A(n33198), .Y(n23544) );
  INVX1 U11819 ( .A(n23544), .Y(n23545) );
  INVX1 U11820 ( .A(n33202), .Y(n23546) );
  INVX1 U11821 ( .A(n23546), .Y(n23547) );
  INVX1 U11822 ( .A(n33205), .Y(n23548) );
  INVX1 U11823 ( .A(n23548), .Y(n23549) );
  BUFX2 U11824 ( .A(n33225), .Y(n23550) );
  BUFX2 U11825 ( .A(n33228), .Y(n23551) );
  INVX1 U11826 ( .A(n33232), .Y(n23552) );
  INVX1 U11827 ( .A(n23552), .Y(n23553) );
  BUFX2 U11828 ( .A(n33236), .Y(n23554) );
  BUFX2 U11829 ( .A(n33256), .Y(n23555) );
  INVX1 U11830 ( .A(n33259), .Y(n23556) );
  INVX1 U11831 ( .A(n23556), .Y(n23557) );
  BUFX2 U11832 ( .A(n33263), .Y(n23558) );
  INVX4 U11833 ( .A(n29439), .Y(n29424) );
  BUFX2 U11834 ( .A(n33266), .Y(n23559) );
  BUFX2 U11835 ( .A(n33286), .Y(n23560) );
  BUFX2 U11836 ( .A(n33289), .Y(n23561) );
  BUFX2 U11837 ( .A(n33293), .Y(n23562) );
  INVX1 U11838 ( .A(n33297), .Y(n23563) );
  INVX1 U11839 ( .A(n23563), .Y(n23564) );
  BUFX2 U11840 ( .A(n33317), .Y(n23565) );
  BUFX2 U11841 ( .A(n33320), .Y(n23566) );
  BUFX2 U11842 ( .A(n33324), .Y(n23567) );
  BUFX2 U11843 ( .A(n33328), .Y(n23568) );
  INVX1 U11844 ( .A(n33348), .Y(n23569) );
  INVX1 U11845 ( .A(n23569), .Y(n23570) );
  BUFX2 U11846 ( .A(n33351), .Y(n23571) );
  BUFX2 U11847 ( .A(n33355), .Y(n23572) );
  INVX1 U11848 ( .A(n33358), .Y(n23573) );
  INVX1 U11849 ( .A(n23573), .Y(n23574) );
  INVX1 U11850 ( .A(n33378), .Y(n23575) );
  INVX1 U11851 ( .A(n23575), .Y(n23576) );
  BUFX2 U11852 ( .A(n33381), .Y(n23577) );
  INVX4 U11853 ( .A(n29393), .Y(n29386) );
  INVX1 U11854 ( .A(n33385), .Y(n23578) );
  INVX1 U11855 ( .A(n23578), .Y(n23579) );
  INVX1 U11856 ( .A(n33388), .Y(n23580) );
  INVX1 U11857 ( .A(n23580), .Y(n23581) );
  BUFX2 U11858 ( .A(n33408), .Y(n23582) );
  INVX4 U11859 ( .A(n29410), .Y(n29408) );
  BUFX2 U11860 ( .A(n33411), .Y(n23583) );
  INVX4 U11861 ( .A(n33885), .Y(n29348) );
  BUFX2 U11862 ( .A(n33415), .Y(n23584) );
  INVX4 U11863 ( .A(n29410), .Y(n29409) );
  BUFX2 U11864 ( .A(n33419), .Y(n23585) );
  INVX4 U11865 ( .A(n29343), .Y(n29349) );
  BUFX2 U11866 ( .A(n33929), .Y(n23586) );
  BUFX2 U11867 ( .A(n34285), .Y(n23587) );
  BUFX2 U11868 ( .A(n34345), .Y(n23588) );
  INVX4 U11869 ( .A(n29411), .Y(n29407) );
  BUFX2 U11870 ( .A(n29635), .Y(n23589) );
  BUFX2 U11871 ( .A(n29695), .Y(n23590) );
  BUFX2 U11872 ( .A(n29705), .Y(n23591) );
  BUFX2 U11873 ( .A(n30043), .Y(n23592) );
  BUFX2 U11874 ( .A(n16209), .Y(n23593) );
  BUFX2 U11875 ( .A(n16128), .Y(n23594) );
  BUFX2 U11876 ( .A(n16051), .Y(n23595) );
  BUFX2 U11877 ( .A(n15977), .Y(n23596) );
  INVX1 U11878 ( .A(n33194), .Y(n23597) );
  INVX1 U11879 ( .A(n23597), .Y(n23598) );
  INVX1 U11880 ( .A(n33296), .Y(n23599) );
  INVX1 U11881 ( .A(n23599), .Y(n23600) );
  INVX1 U11882 ( .A(n34200), .Y(n23601) );
  INVX1 U11883 ( .A(n23601), .Y(n23602) );
  AND2X2 U11884 ( .A(n29068), .B(n2255), .Y(n25523) );
  INVX1 U11885 ( .A(n25523), .Y(n23603) );
  INVX1 U11886 ( .A(n29710), .Y(n23604) );
  INVX1 U11887 ( .A(n23604), .Y(n23605) );
  INVX1 U11888 ( .A(n31056), .Y(n23606) );
  INVX1 U11889 ( .A(n23606), .Y(n23607) );
  INVX1 U11890 ( .A(n34208), .Y(n23608) );
  INVX1 U11891 ( .A(n23608), .Y(n23609) );
  INVX1 U11892 ( .A(n33923), .Y(n23610) );
  INVX4 U11893 ( .A(n23610), .Y(n23611) );
  INVX1 U11894 ( .A(n29563), .Y(n33923) );
  INVX1 U11895 ( .A(n30459), .Y(n23612) );
  INVX2 U11896 ( .A(n23612), .Y(n23613) );
  INVX1 U11897 ( .A(n30120), .Y(n30459) );
  INVX1 U11898 ( .A(n23292), .Y(n23614) );
  INVX1 U11899 ( .A(n32631), .Y(n23615) );
  INVX1 U11900 ( .A(n23615), .Y(n23616) );
  INVX1 U11901 ( .A(n34247), .Y(n25762) );
  INVX1 U11902 ( .A(n30938), .Y(n23618) );
  INVX1 U11903 ( .A(n30940), .Y(n23619) );
  INVX1 U11904 ( .A(n31016), .Y(n23621) );
  INVX1 U11905 ( .A(n31018), .Y(n23622) );
  INVX1 U11906 ( .A(n31583), .Y(n23624) );
  INVX1 U11907 ( .A(n31585), .Y(n23625) );
  AND2X2 U11908 ( .A(n21534), .B(n23940), .Y(n21822) );
  INVX1 U11909 ( .A(n21822), .Y(n23627) );
  AND2X2 U11910 ( .A(n21536), .B(n23943), .Y(n21817) );
  INVX1 U11911 ( .A(n21817), .Y(n23628) );
  OR2X1 U11912 ( .A(n29370), .B(n34159), .Y(n21770) );
  INVX1 U11913 ( .A(n21770), .Y(n23629) );
  AND2X2 U11914 ( .A(n21552), .B(n23998), .Y(n20539) );
  INVX1 U11915 ( .A(n20539), .Y(n23630) );
  AND2X2 U11916 ( .A(n21539), .B(n23903), .Y(n20537) );
  INVX1 U11917 ( .A(n20537), .Y(n23631) );
  AND2X2 U11918 ( .A(n21541), .B(n23945), .Y(n21847) );
  INVX1 U11919 ( .A(n21847), .Y(n23632) );
  INVX1 U11920 ( .A(n23273), .Y(n23633) );
  INVX1 U11921 ( .A(n32475), .Y(n25746) );
  INVX1 U11922 ( .A(n23611), .Y(n23635) );
  INVX1 U11923 ( .A(n30127), .Y(n23636) );
  INVX1 U11924 ( .A(n34189), .Y(n23637) );
  INVX4 U11925 ( .A(n33928), .Y(n30127) );
  OR2X1 U11926 ( .A(n25217), .B(n25218), .Y(n25216) );
  INVX1 U11927 ( .A(n25216), .Y(n23639) );
  OR2X1 U11928 ( .A(n16140), .B(n16139), .Y(n25218) );
  OR2X1 U11929 ( .A(n25220), .B(n25221), .Y(n25219) );
  OR2X1 U11930 ( .A(n16063), .B(n16062), .Y(n25221) );
  AND2X2 U11931 ( .A(n27903), .B(n29189), .Y(n25588) );
  AND2X2 U11932 ( .A(n21546), .B(n23921), .Y(n27143) );
  AND2X1 U11933 ( .A(data_in[4]), .B(data_in[0]), .Y(n31868) );
  AND2X1 U11934 ( .A(n27273), .B(n26708), .Y(n29751) );
  AND2X2 U11935 ( .A(n3209), .B(n32528), .Y(n32906) );
  INVX1 U11936 ( .A(n32906), .Y(n23640) );
  OR2X1 U11937 ( .A(n16122), .B(n34583), .Y(n16093) );
  INVX1 U11938 ( .A(n16093), .Y(n23641) );
  OR2X1 U11939 ( .A(n15971), .B(n34573), .Y(n15942) );
  INVX1 U11940 ( .A(n15942), .Y(n23642) );
  AND2X1 U11941 ( .A(n34603), .B(n29217), .Y(n30480) );
  INVX1 U11942 ( .A(n30480), .Y(n23643) );
  INVX1 U11943 ( .A(n25617), .Y(n23644) );
  INVX1 U11944 ( .A(n25195), .Y(n23645) );
  BUFX2 U11945 ( .A(n29482), .Y(n23646) );
  BUFX2 U11946 ( .A(n29634), .Y(n23647) );
  BUFX2 U11947 ( .A(n30042), .Y(n23648) );
  BUFX2 U11948 ( .A(n30083), .Y(n23649) );
  BUFX2 U11949 ( .A(n30090), .Y(n23650) );
  BUFX2 U11950 ( .A(n30098), .Y(n23651) );
  BUFX2 U11951 ( .A(n30107), .Y(n23652) );
  BUFX2 U11952 ( .A(n30115), .Y(n23653) );
  BUFX2 U11953 ( .A(n30124), .Y(n23654) );
  BUFX2 U11954 ( .A(n30133), .Y(n23655) );
  BUFX2 U11955 ( .A(n30141), .Y(n23656) );
  BUFX2 U11956 ( .A(n30147), .Y(n23657) );
  BUFX2 U11957 ( .A(n30152), .Y(n23658) );
  BUFX2 U11958 ( .A(n30157), .Y(n23659) );
  BUFX2 U11959 ( .A(n30162), .Y(n23660) );
  BUFX2 U11960 ( .A(n30167), .Y(n23661) );
  BUFX2 U11961 ( .A(n30172), .Y(n23662) );
  BUFX2 U11962 ( .A(n30177), .Y(n23663) );
  BUFX2 U11963 ( .A(n30183), .Y(n23664) );
  BUFX2 U11964 ( .A(n30193), .Y(n23665) );
  BUFX2 U11965 ( .A(n30198), .Y(n23666) );
  BUFX2 U11966 ( .A(n30203), .Y(n23667) );
  BUFX2 U11967 ( .A(n30208), .Y(n23668) );
  BUFX2 U11968 ( .A(n30213), .Y(n23669) );
  BUFX2 U11969 ( .A(n30218), .Y(n23670) );
  BUFX2 U11970 ( .A(n30223), .Y(n23671) );
  BUFX2 U11971 ( .A(n30232), .Y(n23672) );
  BUFX2 U11972 ( .A(n30241), .Y(n23673) );
  BUFX2 U11973 ( .A(n30246), .Y(n23674) );
  BUFX2 U11974 ( .A(n30251), .Y(n23675) );
  BUFX2 U11975 ( .A(n30256), .Y(n23676) );
  BUFX2 U11976 ( .A(n30261), .Y(n23677) );
  BUFX2 U11977 ( .A(n30266), .Y(n23678) );
  BUFX2 U11978 ( .A(n30270), .Y(n23679) );
  BUFX2 U11979 ( .A(n30278), .Y(n23680) );
  BUFX2 U11980 ( .A(n30287), .Y(n23681) );
  BUFX2 U11981 ( .A(n30292), .Y(n23682) );
  BUFX2 U11982 ( .A(n30297), .Y(n23683) );
  BUFX2 U11983 ( .A(n30302), .Y(n23684) );
  BUFX2 U11984 ( .A(n30307), .Y(n23685) );
  BUFX2 U11985 ( .A(n30312), .Y(n23686) );
  BUFX2 U11986 ( .A(n30317), .Y(n23687) );
  BUFX2 U11987 ( .A(n30325), .Y(n23688) );
  BUFX2 U11988 ( .A(n30333), .Y(n23689) );
  BUFX2 U11989 ( .A(n30338), .Y(n23690) );
  BUFX2 U11990 ( .A(n30343), .Y(n23691) );
  BUFX2 U11991 ( .A(n30347), .Y(n23692) );
  BUFX2 U11992 ( .A(n30352), .Y(n23693) );
  BUFX2 U11993 ( .A(n30357), .Y(n23694) );
  BUFX2 U11994 ( .A(n30362), .Y(n23695) );
  BUFX2 U11995 ( .A(n30369), .Y(n23696) );
  BUFX2 U11996 ( .A(n30378), .Y(n23697) );
  BUFX2 U11997 ( .A(n30383), .Y(n23698) );
  BUFX2 U11998 ( .A(n30387), .Y(n23699) );
  BUFX2 U11999 ( .A(n30392), .Y(n23700) );
  BUFX2 U12000 ( .A(n30397), .Y(n23701) );
  BUFX2 U12001 ( .A(n30402), .Y(n23702) );
  BUFX2 U12002 ( .A(n30407), .Y(n23703) );
  BUFX2 U12003 ( .A(n30416), .Y(n23704) );
  BUFX2 U12004 ( .A(n30424), .Y(n23705) );
  BUFX2 U12005 ( .A(n30430), .Y(n23706) );
  BUFX2 U12006 ( .A(n30438), .Y(n23707) );
  BUFX2 U12007 ( .A(n30447), .Y(n23708) );
  BUFX2 U12008 ( .A(n30455), .Y(n23709) );
  BUFX2 U12009 ( .A(n30462), .Y(n23710) );
  BUFX2 U12010 ( .A(n30469), .Y(n23711) );
  BUFX2 U12011 ( .A(n33197), .Y(n23712) );
  BUFX2 U12012 ( .A(n33204), .Y(n23713) );
  BUFX2 U12013 ( .A(n33224), .Y(n23714) );
  BUFX2 U12014 ( .A(n33227), .Y(n23715) );
  BUFX2 U12015 ( .A(n33235), .Y(n23716) );
  BUFX2 U12016 ( .A(n33255), .Y(n23717) );
  BUFX2 U12017 ( .A(n33258), .Y(n23718) );
  INVX4 U12018 ( .A(n29402), .Y(n29398) );
  BUFX2 U12019 ( .A(n33265), .Y(n23719) );
  BUFX2 U12020 ( .A(n33285), .Y(n23720) );
  BUFX2 U12021 ( .A(n33288), .Y(n23721) );
  BUFX2 U12022 ( .A(n33292), .Y(n23722) );
  BUFX2 U12023 ( .A(n33316), .Y(n23723) );
  BUFX2 U12024 ( .A(n33319), .Y(n23724) );
  BUFX2 U12025 ( .A(n33323), .Y(n23725) );
  INVX4 U12026 ( .A(n29354), .Y(n29359) );
  BUFX2 U12027 ( .A(n33327), .Y(n23726) );
  BUFX2 U12028 ( .A(n33347), .Y(n23727) );
  INVX4 U12029 ( .A(n34219), .Y(n29361) );
  BUFX2 U12030 ( .A(n33350), .Y(n23728) );
  BUFX2 U12031 ( .A(n33354), .Y(n23729) );
  BUFX2 U12032 ( .A(n33357), .Y(n23730) );
  BUFX2 U12033 ( .A(n33377), .Y(n23731) );
  INVX4 U12034 ( .A(n34219), .Y(n29362) );
  BUFX2 U12035 ( .A(n33380), .Y(n23732) );
  BUFX2 U12036 ( .A(n33387), .Y(n23733) );
  BUFX2 U12037 ( .A(n33407), .Y(n23734) );
  BUFX2 U12038 ( .A(n33410), .Y(n23735) );
  BUFX2 U12039 ( .A(n33414), .Y(n23736) );
  BUFX2 U12040 ( .A(n33418), .Y(n23737) );
  INVX4 U12041 ( .A(n29402), .Y(n29396) );
  BUFX2 U12042 ( .A(n34284), .Y(n23738) );
  INVX4 U12043 ( .A(n29402), .Y(n29397) );
  BUFX2 U12044 ( .A(n34344), .Y(n23739) );
  BUFX2 U12045 ( .A(n16210), .Y(n23740) );
  BUFX2 U12046 ( .A(n16129), .Y(n23741) );
  BUFX2 U12047 ( .A(n16052), .Y(n23742) );
  BUFX2 U12048 ( .A(n15978), .Y(n23743) );
  AND2X2 U12049 ( .A(n27281), .B(net96596), .Y(n25521) );
  INVX1 U12050 ( .A(n25521), .Y(n23744) );
  INVX1 U12051 ( .A(n29711), .Y(n23745) );
  OR2X2 U12052 ( .A(n23605), .B(n22130), .Y(n29711) );
  AND2X2 U12053 ( .A(n11684), .B(net96578), .Y(n34288) );
  INVX1 U12054 ( .A(n34288), .Y(n23746) );
  INVX1 U12055 ( .A(n29515), .Y(n23747) );
  INVX1 U12056 ( .A(n23747), .Y(n23748) );
  BUFX2 U12057 ( .A(n29761), .Y(n23749) );
  BUFX2 U12058 ( .A(n29770), .Y(n23750) );
  BUFX2 U12059 ( .A(n29778), .Y(n23751) );
  BUFX2 U12060 ( .A(n29786), .Y(n23752) );
  BUFX2 U12061 ( .A(n29795), .Y(n23753) );
  BUFX2 U12062 ( .A(n29804), .Y(n23754) );
  BUFX2 U12063 ( .A(n29816), .Y(n23755) );
  BUFX2 U12064 ( .A(n29826), .Y(n23756) );
  BUFX2 U12065 ( .A(n29837), .Y(n23757) );
  BUFX2 U12066 ( .A(n29847), .Y(n23758) );
  BUFX2 U12067 ( .A(n29855), .Y(n23759) );
  BUFX2 U12068 ( .A(n29863), .Y(n23760) );
  BUFX2 U12069 ( .A(n29872), .Y(n23761) );
  BUFX2 U12070 ( .A(n29900), .Y(n23762) );
  BUFX2 U12071 ( .A(n29910), .Y(n23763) );
  BUFX2 U12072 ( .A(n29920), .Y(n23764) );
  BUFX2 U12073 ( .A(n29931), .Y(n23765) );
  BUFX2 U12074 ( .A(n29941), .Y(n23766) );
  BUFX2 U12075 ( .A(n29954), .Y(n23767) );
  BUFX2 U12076 ( .A(n29964), .Y(n23768) );
  BUFX2 U12077 ( .A(n29976), .Y(n23769) );
  BUFX2 U12078 ( .A(n29987), .Y(n23770) );
  BUFX2 U12079 ( .A(n29999), .Y(n23771) );
  BUFX2 U12080 ( .A(n30010), .Y(n23772) );
  BUFX2 U12081 ( .A(n30020), .Y(n23773) );
  BUFX2 U12082 ( .A(n32628), .Y(n23774) );
  INVX4 U12083 ( .A(n25454), .Y(n33369) );
  BUFX2 U12084 ( .A(n32635), .Y(n23775) );
  INVX4 U12085 ( .A(n25430), .Y(n33295) );
  BUFX2 U12086 ( .A(n32713), .Y(n23776) );
  BUFX2 U12087 ( .A(n32723), .Y(n23777) );
  BUFX2 U12088 ( .A(n32908), .Y(n23778) );
  INVX4 U12089 ( .A(n21160), .Y(n33399) );
  BUFX2 U12090 ( .A(n32930), .Y(n23779) );
  INVX4 U12091 ( .A(n25425), .Y(n33508) );
  INVX8 U12092 ( .A(n25427), .Y(n33485) );
  BUFX2 U12093 ( .A(n32951), .Y(n23780) );
  INVX4 U12094 ( .A(n27022), .Y(n33639) );
  BUFX2 U12095 ( .A(n33017), .Y(n23781) );
  INVX4 U12096 ( .A(n25352), .Y(n33430) );
  BUFX2 U12097 ( .A(n33020), .Y(n23782) );
  INVX4 U12098 ( .A(n25354), .Y(n33339) );
  BUFX2 U12099 ( .A(n33037), .Y(n23783) );
  INVX4 U12100 ( .A(n25423), .Y(n33587) );
  INVX4 U12101 ( .A(n25402), .Y(n33551) );
  BUFX2 U12102 ( .A(n33039), .Y(n23784) );
  BUFX2 U12103 ( .A(n29630), .Y(n23785) );
  BUFX2 U12104 ( .A(n29684), .Y(n23786) );
  BUFX2 U12105 ( .A(n29737), .Y(n23787) );
  BUFX2 U12106 ( .A(n29739), .Y(n23788) );
  BUFX2 U12107 ( .A(n29749), .Y(n23789) );
  BUFX2 U12108 ( .A(n29762), .Y(n23790) );
  BUFX2 U12109 ( .A(n29771), .Y(n23791) );
  BUFX2 U12110 ( .A(n29779), .Y(n23792) );
  BUFX2 U12111 ( .A(n29787), .Y(n23793) );
  BUFX2 U12112 ( .A(n29796), .Y(n23794) );
  BUFX2 U12113 ( .A(n29805), .Y(n23795) );
  BUFX2 U12114 ( .A(n29817), .Y(n23796) );
  BUFX2 U12115 ( .A(n29827), .Y(n23797) );
  BUFX2 U12116 ( .A(n29838), .Y(n23798) );
  BUFX2 U12117 ( .A(n29848), .Y(n23799) );
  BUFX2 U12118 ( .A(n29856), .Y(n23800) );
  BUFX2 U12119 ( .A(n29864), .Y(n23801) );
  BUFX2 U12120 ( .A(n29873), .Y(n23802) );
  BUFX2 U12121 ( .A(n29880), .Y(n23803) );
  BUFX2 U12122 ( .A(n29890), .Y(n23804) );
  BUFX2 U12123 ( .A(n29901), .Y(n23805) );
  BUFX2 U12124 ( .A(n29911), .Y(n23806) );
  BUFX2 U12125 ( .A(n29921), .Y(n23807) );
  BUFX2 U12126 ( .A(n29932), .Y(n23808) );
  BUFX2 U12127 ( .A(n29942), .Y(n23809) );
  BUFX2 U12128 ( .A(n29955), .Y(n23810) );
  BUFX2 U12129 ( .A(n29965), .Y(n23811) );
  BUFX2 U12130 ( .A(n29977), .Y(n23812) );
  BUFX2 U12131 ( .A(n29988), .Y(n23813) );
  BUFX2 U12132 ( .A(n30000), .Y(n23814) );
  BUFX2 U12133 ( .A(n30011), .Y(n23815) );
  BUFX2 U12134 ( .A(n30022), .Y(n23816) );
  BUFX2 U12135 ( .A(n30034), .Y(n23817) );
  BUFX2 U12136 ( .A(n30081), .Y(n23818) );
  BUFX2 U12137 ( .A(n30088), .Y(n23819) );
  BUFX2 U12138 ( .A(n30096), .Y(n23820) );
  BUFX2 U12139 ( .A(n30105), .Y(n23821) );
  BUFX2 U12140 ( .A(n30113), .Y(n23822) );
  BUFX2 U12141 ( .A(n30122), .Y(n23823) );
  BUFX2 U12142 ( .A(n30131), .Y(n23824) );
  BUFX2 U12143 ( .A(n30139), .Y(n23825) );
  BUFX2 U12144 ( .A(n30145), .Y(n23826) );
  BUFX2 U12145 ( .A(n30150), .Y(n23827) );
  BUFX2 U12146 ( .A(n30155), .Y(n23828) );
  BUFX2 U12147 ( .A(n30160), .Y(n23829) );
  BUFX2 U12148 ( .A(n30165), .Y(n23830) );
  BUFX2 U12149 ( .A(n30170), .Y(n23831) );
  BUFX2 U12150 ( .A(n30175), .Y(n23832) );
  BUFX2 U12151 ( .A(n30181), .Y(n23833) );
  BUFX2 U12152 ( .A(n30191), .Y(n23834) );
  BUFX2 U12153 ( .A(n30196), .Y(n23835) );
  BUFX2 U12154 ( .A(n30201), .Y(n23836) );
  BUFX2 U12155 ( .A(n30206), .Y(n23837) );
  BUFX2 U12156 ( .A(n30211), .Y(n23838) );
  BUFX2 U12157 ( .A(n30216), .Y(n23839) );
  BUFX2 U12158 ( .A(n30221), .Y(n23840) );
  BUFX2 U12159 ( .A(n30230), .Y(n23841) );
  BUFX2 U12160 ( .A(n30239), .Y(n23842) );
  BUFX2 U12161 ( .A(n30244), .Y(n23843) );
  BUFX2 U12162 ( .A(n30249), .Y(n23844) );
  BUFX2 U12163 ( .A(n30254), .Y(n23845) );
  BUFX2 U12164 ( .A(n30259), .Y(n23846) );
  BUFX2 U12165 ( .A(n30264), .Y(n23847) );
  BUFX2 U12166 ( .A(n30268), .Y(n23848) );
  BUFX2 U12167 ( .A(n30276), .Y(n23849) );
  BUFX2 U12168 ( .A(n30285), .Y(n23850) );
  BUFX2 U12169 ( .A(n30290), .Y(n23851) );
  BUFX2 U12170 ( .A(n30295), .Y(n23852) );
  BUFX2 U12171 ( .A(n30300), .Y(n23853) );
  BUFX2 U12172 ( .A(n30305), .Y(n23854) );
  BUFX2 U12173 ( .A(n30310), .Y(n23855) );
  BUFX2 U12174 ( .A(n30315), .Y(n23856) );
  BUFX2 U12175 ( .A(n30323), .Y(n23857) );
  BUFX2 U12176 ( .A(n30331), .Y(n23858) );
  BUFX2 U12177 ( .A(n30336), .Y(n23859) );
  BUFX2 U12178 ( .A(n30341), .Y(n23860) );
  BUFX2 U12179 ( .A(n30345), .Y(n23861) );
  BUFX2 U12180 ( .A(n30350), .Y(n23862) );
  BUFX2 U12181 ( .A(n30355), .Y(n23863) );
  BUFX2 U12182 ( .A(n30360), .Y(n23864) );
  BUFX2 U12183 ( .A(n30367), .Y(n23865) );
  BUFX2 U12184 ( .A(n30376), .Y(n23866) );
  BUFX2 U12185 ( .A(n30381), .Y(n23867) );
  BUFX2 U12186 ( .A(n30385), .Y(n23868) );
  BUFX2 U12187 ( .A(n30390), .Y(n23869) );
  BUFX2 U12188 ( .A(n30395), .Y(n23870) );
  BUFX2 U12189 ( .A(n30400), .Y(n23871) );
  BUFX2 U12190 ( .A(n30405), .Y(n23872) );
  BUFX2 U12191 ( .A(n30414), .Y(n23873) );
  BUFX2 U12192 ( .A(n30422), .Y(n23874) );
  BUFX2 U12193 ( .A(n30428), .Y(n23875) );
  BUFX2 U12194 ( .A(n30436), .Y(n23876) );
  BUFX2 U12195 ( .A(n30445), .Y(n23877) );
  BUFX2 U12196 ( .A(n30453), .Y(n23878) );
  BUFX2 U12197 ( .A(n30460), .Y(n23879) );
  BUFX2 U12198 ( .A(n30467), .Y(n23880) );
  BUFX2 U12199 ( .A(n33160), .Y(n23881) );
  BUFX2 U12200 ( .A(n33372), .Y(n23882) );
  INVX4 U12201 ( .A(n29401), .Y(n29400) );
  BUFX2 U12202 ( .A(n34223), .Y(n23883) );
  BUFX2 U12203 ( .A(n16194), .Y(n23884) );
  BUFX2 U12204 ( .A(n16113), .Y(n23885) );
  BUFX2 U12205 ( .A(n16036), .Y(n23886) );
  BUFX2 U12206 ( .A(n15962), .Y(n23887) );
  INVX1 U12207 ( .A(n25195), .Y(n23888) );
  AND2X2 U12208 ( .A(n34385), .B(n33069), .Y(n25697) );
  AND2X1 U12209 ( .A(n30021), .B(n24976), .Y(n29896) );
  INVX1 U12210 ( .A(n29896), .Y(n23889) );
  AND2X2 U12211 ( .A(n29440), .B(n32463), .Y(n30481) );
  INVX1 U12212 ( .A(n30481), .Y(n23890) );
  AND2X1 U12213 ( .A(n16183), .B(n25214), .Y(n16182) );
  INVX1 U12214 ( .A(n16182), .Y(n23891) );
  AND2X1 U12215 ( .A(n16109), .B(n25197), .Y(n16108) );
  INVX1 U12216 ( .A(n16108), .Y(n23892) );
  AND2X1 U12217 ( .A(n16102), .B(n23639), .Y(n16101) );
  INVX1 U12218 ( .A(n16101), .Y(n23893) );
  AND2X1 U12219 ( .A(n16025), .B(n34596), .Y(n16024) );
  INVX1 U12220 ( .A(n16024), .Y(n23894) );
  AND2X1 U12221 ( .A(n15958), .B(n25199), .Y(n15957) );
  INVX1 U12222 ( .A(n15957), .Y(n23895) );
  AND2X1 U12223 ( .A(n15951), .B(n34576), .Y(n15950) );
  INVX1 U12224 ( .A(n15950), .Y(n23896) );
  INVX1 U12225 ( .A(n32171), .Y(n23897) );
  INVX1 U12226 ( .A(n23897), .Y(n23898) );
  INVX1 U12227 ( .A(n32176), .Y(n23899) );
  INVX1 U12228 ( .A(n23899), .Y(n23900) );
  BUFX2 U12229 ( .A(n32181), .Y(n23901) );
  AND2X2 U12230 ( .A(n34174), .B(n27304), .Y(n27263) );
  BUFX2 U12231 ( .A(n34183), .Y(n23902) );
  BUFX2 U12232 ( .A(n34216), .Y(n23903) );
  BUFX2 U12233 ( .A(n15900), .Y(n23904) );
  BUFX2 U12234 ( .A(n29878), .Y(n23905) );
  BUFX2 U12235 ( .A(n29909), .Y(n23906) );
  BUFX2 U12236 ( .A(n29919), .Y(n23907) );
  BUFX2 U12237 ( .A(n29930), .Y(n23908) );
  BUFX2 U12238 ( .A(n29940), .Y(n23909) );
  BUFX2 U12239 ( .A(n29953), .Y(n23910) );
  BUFX2 U12240 ( .A(n29963), .Y(n23911) );
  BUFX2 U12241 ( .A(n29975), .Y(n23912) );
  BUFX2 U12242 ( .A(n29986), .Y(n23913) );
  BUFX2 U12243 ( .A(n29998), .Y(n23914) );
  BUFX2 U12244 ( .A(n30009), .Y(n23915) );
  BUFX2 U12245 ( .A(n30019), .Y(n23916) );
  BUFX2 U12246 ( .A(n30032), .Y(n23917) );
  AND2X2 U12247 ( .A(n29071), .B(n29185), .Y(n25526) );
  INVX1 U12248 ( .A(n25526), .Y(n23918) );
  AND2X2 U12249 ( .A(n27178), .B(n20961), .Y(n26063) );
  INVX1 U12250 ( .A(n26063), .Y(n23919) );
  AND2X2 U12251 ( .A(n3179), .B(n26518), .Y(n27044) );
  INVX1 U12252 ( .A(n27044), .Y(n23920) );
  AND2X2 U12253 ( .A(n33762), .B(n3139), .Y(n27145) );
  INVX1 U12254 ( .A(n27145), .Y(n23921) );
  INVX1 U12255 ( .A(n29718), .Y(n23922) );
  OR2X2 U12256 ( .A(n22113), .B(n22134), .Y(n29718) );
  AND2X2 U12257 ( .A(n3244), .B(n33326), .Y(n32633) );
  INVX1 U12258 ( .A(n32633), .Y(n23923) );
  INVX4 U12259 ( .A(n25428), .Y(n33326) );
  AND2X2 U12260 ( .A(n11682), .B(net96576), .Y(n33935) );
  INVX1 U12261 ( .A(n33935), .Y(n23924) );
  AND2X2 U12262 ( .A(n11681), .B(net96576), .Y(n33937) );
  INVX1 U12263 ( .A(n33937), .Y(n23925) );
  AND2X2 U12264 ( .A(n11679), .B(net96576), .Y(n33941) );
  INVX1 U12265 ( .A(n33941), .Y(n23926) );
  AND2X2 U12266 ( .A(n11678), .B(net96576), .Y(n33943) );
  INVX1 U12267 ( .A(n33943), .Y(n23927) );
  AND2X2 U12268 ( .A(n11677), .B(net96576), .Y(n33945) );
  INVX1 U12269 ( .A(n33945), .Y(n23928) );
  AND2X2 U12270 ( .A(n11674), .B(net96576), .Y(n33951) );
  INVX1 U12271 ( .A(n33951), .Y(n23929) );
  AND2X2 U12272 ( .A(n11673), .B(net96578), .Y(n33953) );
  INVX1 U12273 ( .A(n33953), .Y(n23930) );
  AND2X2 U12274 ( .A(n11670), .B(net96576), .Y(n33957) );
  INVX1 U12275 ( .A(n33957), .Y(n23931) );
  AND2X2 U12276 ( .A(n11669), .B(net96576), .Y(n33959) );
  INVX1 U12277 ( .A(n33959), .Y(n23932) );
  AND2X2 U12278 ( .A(n11668), .B(net96576), .Y(n33961) );
  INVX1 U12279 ( .A(n33961), .Y(n23933) );
  AND2X2 U12280 ( .A(n11667), .B(net96576), .Y(n33963) );
  INVX1 U12281 ( .A(n33963), .Y(n23934) );
  AND2X2 U12282 ( .A(n11665), .B(net96576), .Y(n33967) );
  INVX1 U12283 ( .A(n33967), .Y(n23935) );
  AND2X2 U12284 ( .A(n11664), .B(net96578), .Y(n33969) );
  INVX1 U12285 ( .A(n33969), .Y(n23936) );
  AND2X2 U12286 ( .A(n11663), .B(net96576), .Y(n33971) );
  INVX1 U12287 ( .A(n33971), .Y(n23937) );
  AND2X2 U12288 ( .A(n11662), .B(net96578), .Y(n33972) );
  INVX1 U12289 ( .A(n33972), .Y(n23938) );
  AND2X2 U12290 ( .A(n11661), .B(net96578), .Y(n33974) );
  INVX1 U12291 ( .A(n33974), .Y(n23939) );
  AND2X2 U12292 ( .A(n11660), .B(net96578), .Y(n33976) );
  INVX1 U12293 ( .A(n33976), .Y(n23940) );
  AND2X2 U12294 ( .A(n11659), .B(net96578), .Y(n33978) );
  INVX1 U12295 ( .A(n33978), .Y(n23941) );
  AND2X2 U12296 ( .A(n11657), .B(net96578), .Y(n33982) );
  INVX1 U12297 ( .A(n33982), .Y(n23942) );
  AND2X2 U12298 ( .A(n11655), .B(net96578), .Y(n33986) );
  INVX1 U12299 ( .A(n33986), .Y(n23943) );
  AND2X2 U12300 ( .A(n11683), .B(net96578), .Y(n33988) );
  INVX1 U12301 ( .A(n33988), .Y(n23944) );
  AND2X2 U12302 ( .A(n11685), .B(net96578), .Y(n34347) );
  INVX1 U12303 ( .A(n34347), .Y(n23945) );
  BUFX2 U12304 ( .A(n29632), .Y(n23946) );
  BUFX2 U12305 ( .A(n31895), .Y(n23947) );
  INVX1 U12306 ( .A(n32162), .Y(n23948) );
  INVX1 U12307 ( .A(n23948), .Y(n23949) );
  INVX1 U12308 ( .A(n32167), .Y(n23950) );
  INVX1 U12309 ( .A(n23950), .Y(n23951) );
  INVX1 U12310 ( .A(n32172), .Y(n23952) );
  INVX1 U12311 ( .A(n23952), .Y(n23953) );
  INVX1 U12312 ( .A(n32177), .Y(n23954) );
  INVX1 U12313 ( .A(n23954), .Y(n23955) );
  INVX1 U12314 ( .A(n32182), .Y(n23956) );
  INVX1 U12315 ( .A(n23956), .Y(n23957) );
  INVX1 U12316 ( .A(n32634), .Y(n23958) );
  INVX1 U12317 ( .A(n23958), .Y(n23959) );
  BUFX2 U12318 ( .A(n33433), .Y(n23960) );
  BUFX2 U12319 ( .A(n33446), .Y(n23961) );
  BUFX2 U12320 ( .A(n33451), .Y(n23962) );
  BUFX2 U12321 ( .A(n33468), .Y(n23963) );
  BUFX2 U12322 ( .A(n33474), .Y(n23964) );
  BUFX2 U12323 ( .A(n33491), .Y(n23965) );
  BUFX2 U12324 ( .A(n33497), .Y(n23966) );
  BUFX2 U12325 ( .A(n33514), .Y(n23967) );
  BUFX2 U12326 ( .A(n33520), .Y(n23968) );
  BUFX2 U12327 ( .A(n33570), .Y(n23969) );
  BUFX2 U12328 ( .A(n33576), .Y(n23970) );
  BUFX2 U12329 ( .A(n33593), .Y(n23971) );
  BUFX2 U12330 ( .A(n33598), .Y(n23972) );
  BUFX2 U12331 ( .A(n33615), .Y(n23973) );
  BUFX2 U12332 ( .A(n33620), .Y(n23974) );
  BUFX2 U12333 ( .A(n33636), .Y(n23975) );
  BUFX2 U12334 ( .A(n33642), .Y(n23976) );
  BUFX2 U12335 ( .A(n33659), .Y(n23977) );
  BUFX2 U12336 ( .A(n33664), .Y(n23978) );
  BUFX2 U12337 ( .A(n33680), .Y(n23979) );
  BUFX2 U12338 ( .A(n33685), .Y(n23980) );
  BUFX2 U12339 ( .A(n33707), .Y(n23981) );
  BUFX2 U12340 ( .A(n33724), .Y(n23982) );
  BUFX2 U12341 ( .A(n33729), .Y(n23983) );
  BUFX2 U12342 ( .A(n33745), .Y(n23984) );
  BUFX2 U12343 ( .A(n33768), .Y(n23985) );
  BUFX2 U12344 ( .A(n33773), .Y(n23986) );
  BUFX2 U12345 ( .A(n33790), .Y(n23987) );
  BUFX2 U12346 ( .A(n33795), .Y(n23988) );
  BUFX2 U12347 ( .A(n33835), .Y(n23989) );
  BUFX2 U12348 ( .A(n33840), .Y(n23990) );
  BUFX2 U12349 ( .A(n33858), .Y(n23991) );
  BUFX2 U12350 ( .A(n33864), .Y(n23992) );
  BUFX2 U12351 ( .A(n33881), .Y(n23993) );
  BUFX2 U12352 ( .A(n33924), .Y(n23994) );
  AND2X2 U12353 ( .A(n11656), .B(net96578), .Y(n33984) );
  INVX1 U12354 ( .A(n33984), .Y(n23995) );
  AND2X2 U12355 ( .A(n11654), .B(net96578), .Y(n33990) );
  INVX1 U12356 ( .A(n33990), .Y(n23996) );
  BUFX2 U12357 ( .A(n34190), .Y(n23997) );
  BUFX2 U12358 ( .A(n34204), .Y(n23998) );
  BUFX2 U12359 ( .A(n33702), .Y(n23999) );
  BUFX2 U12360 ( .A(n33751), .Y(n24000) );
  BUFX2 U12361 ( .A(n33812), .Y(n24001) );
  BUFX2 U12362 ( .A(n33818), .Y(n24002) );
  BUFX2 U12363 ( .A(n33888), .Y(n24003) );
  INVX1 U12364 ( .A(n25469), .Y(n24004) );
  INVX1 U12365 ( .A(n25471), .Y(n24005) );
  AND2X2 U12366 ( .A(n29052), .B(n29476), .Y(n25470) );
  INVX1 U12367 ( .A(n25470), .Y(n24006) );
  AND2X2 U12368 ( .A(n29083), .B(n29476), .Y(n25522) );
  INVX1 U12369 ( .A(n25522), .Y(n24007) );
  AND2X2 U12370 ( .A(n29074), .B(n29465), .Y(n25525) );
  INVX1 U12371 ( .A(n25525), .Y(n24008) );
  AND2X2 U12372 ( .A(n11680), .B(net96576), .Y(n33939) );
  INVX1 U12373 ( .A(n33939), .Y(n24009) );
  AND2X2 U12374 ( .A(n11676), .B(net96576), .Y(n33947) );
  INVX1 U12375 ( .A(n33947), .Y(n24010) );
  AND2X2 U12376 ( .A(n11675), .B(net96576), .Y(n33949) );
  INVX1 U12377 ( .A(n33949), .Y(n24011) );
  AND2X2 U12378 ( .A(n11671), .B(net96576), .Y(n33955) );
  INVX1 U12379 ( .A(n33955), .Y(n24012) );
  AND2X2 U12380 ( .A(n11666), .B(net96576), .Y(n33965) );
  INVX1 U12381 ( .A(n33965), .Y(n24013) );
  INVX1 U12382 ( .A(n32823), .Y(n24014) );
  INVX1 U12383 ( .A(n24014), .Y(n24015) );
  BUFX2 U12384 ( .A(n16073), .Y(n24016) );
  INVX1 U12385 ( .A(n30484), .Y(n24017) );
  OR2X1 U12386 ( .A(n16075), .B(n15921), .Y(n16074) );
  INVX1 U12387 ( .A(n16074), .Y(n24018) );
  AND2X2 U12388 ( .A(n23543), .B(n23598), .Y(n27292) );
  AND2X2 U12389 ( .A(n23547), .B(n21548), .Y(n27293) );
  AND2X2 U12390 ( .A(n23550), .B(n23714), .Y(n27284) );
  AND2X2 U12391 ( .A(n23553), .B(n21549), .Y(n27287) );
  AND2X2 U12392 ( .A(n23555), .B(n23717), .Y(n27277) );
  AND2X2 U12393 ( .A(n23558), .B(n23430), .Y(n27278) );
  AND2X2 U12394 ( .A(n23560), .B(n23720), .Y(n27279) );
  AND2X2 U12395 ( .A(n23562), .B(n23722), .Y(n27280) );
  AND2X2 U12396 ( .A(n23565), .B(n23723), .Y(n27285) );
  AND2X2 U12397 ( .A(n23567), .B(n23725), .Y(n27288) );
  AND2X2 U12398 ( .A(n23570), .B(n23727), .Y(n27286) );
  AND2X2 U12399 ( .A(n23572), .B(n23729), .Y(n27289) );
  AND2X2 U12400 ( .A(n23576), .B(n23731), .Y(n27290) );
  AND2X2 U12401 ( .A(n23582), .B(n23734), .Y(n27282) );
  AND2X2 U12402 ( .A(n23584), .B(n23736), .Y(n27291) );
  AND2X2 U12403 ( .A(n23588), .B(n23739), .Y(n27283) );
  BUFX2 U12404 ( .A(n16081), .Y(n24019) );
  BUFX2 U12405 ( .A(n15928), .Y(n24020) );
  BUFX2 U12406 ( .A(n16151), .Y(n24021) );
  BUFX2 U12407 ( .A(n16150), .Y(n24022) );
  BUFX2 U12408 ( .A(n16148), .Y(n24023) );
  BUFX2 U12409 ( .A(n16079), .Y(n24024) );
  BUFX2 U12410 ( .A(n16077), .Y(n24025) );
  BUFX2 U12411 ( .A(n16076), .Y(n24026) );
  BUFX2 U12412 ( .A(n16000), .Y(n24027) );
  BUFX2 U12413 ( .A(n15999), .Y(n24028) );
  BUFX2 U12414 ( .A(n15997), .Y(n24029) );
  BUFX2 U12415 ( .A(n15926), .Y(n24030) );
  BUFX2 U12416 ( .A(n15924), .Y(n24031) );
  BUFX2 U12417 ( .A(n15922), .Y(n24032) );
  AND2X2 U12418 ( .A(n23443), .B(n25210), .Y(n30053) );
  INVX1 U12419 ( .A(n30053), .Y(n24033) );
  AND2X2 U12420 ( .A(n23118), .B(n23006), .Y(n30797) );
  INVX1 U12421 ( .A(n30797), .Y(n24034) );
  AND2X2 U12422 ( .A(n23133), .B(n25171), .Y(n30897) );
  INVX1 U12423 ( .A(n30897), .Y(n24035) );
  AND2X2 U12424 ( .A(n23119), .B(n23011), .Y(n30918) );
  INVX1 U12425 ( .A(n30918), .Y(n24036) );
  AND2X2 U12426 ( .A(n23120), .B(n25173), .Y(n30958) );
  INVX1 U12427 ( .A(n30958), .Y(n24037) );
  AND2X2 U12428 ( .A(n23122), .B(n25174), .Y(n31133) );
  INVX1 U12429 ( .A(n31133), .Y(n24038) );
  AND2X2 U12430 ( .A(n23081), .B(n25178), .Y(n31288) );
  INVX1 U12431 ( .A(n31288), .Y(n24039) );
  AND2X2 U12432 ( .A(n23083), .B(n23035), .Y(n31307) );
  INVX1 U12433 ( .A(n31307), .Y(n24040) );
  AND2X2 U12434 ( .A(n23123), .B(n25179), .Y(n31344) );
  INVX1 U12435 ( .A(n31344), .Y(n24041) );
  AND2X2 U12436 ( .A(n23125), .B(n23038), .Y(n31364) );
  INVX1 U12437 ( .A(n31364), .Y(n24042) );
  AND2X2 U12438 ( .A(n25180), .B(n23135), .Y(n31384) );
  INVX1 U12439 ( .A(n31384), .Y(n24043) );
  AND2X2 U12440 ( .A(n23137), .B(n25181), .Y(n31464) );
  INVX1 U12441 ( .A(n31464), .Y(n24044) );
  AND2X2 U12442 ( .A(n23129), .B(n23061), .Y(n31793) );
  INVX1 U12443 ( .A(n31793), .Y(n24045) );
  AND2X2 U12444 ( .A(n23131), .B(n23065), .Y(n31832) );
  INVX1 U12445 ( .A(n31832), .Y(n24046) );
  BUFX2 U12446 ( .A(n30649), .Y(n24047) );
  INVX1 U12447 ( .A(n30840), .Y(n24048) );
  INVX1 U12448 ( .A(n24048), .Y(n24049) );
  INVX1 U12449 ( .A(n30900), .Y(n24050) );
  INVX1 U12450 ( .A(n24050), .Y(n24051) );
  INVX1 U12451 ( .A(n30961), .Y(n24052) );
  INVX1 U12452 ( .A(n24052), .Y(n24053) );
  INVX1 U12453 ( .A(n31005), .Y(n24054) );
  INVX1 U12454 ( .A(n24054), .Y(n24055) );
  INVX1 U12455 ( .A(n31043), .Y(n24056) );
  INVX1 U12456 ( .A(n24056), .Y(n24057) );
  INVX1 U12457 ( .A(n31136), .Y(n24058) );
  INVX1 U12458 ( .A(n24058), .Y(n24059) );
  INVX1 U12459 ( .A(n31161), .Y(n24060) );
  INVX1 U12460 ( .A(n24060), .Y(n24061) );
  INVX1 U12461 ( .A(n31174), .Y(n24062) );
  INVX1 U12462 ( .A(n24062), .Y(n24063) );
  INVX1 U12463 ( .A(n31239), .Y(n24064) );
  INVX1 U12464 ( .A(n24064), .Y(n24065) );
  INVX1 U12465 ( .A(n31279), .Y(n24066) );
  INVX1 U12466 ( .A(n24066), .Y(n24067) );
  INVX1 U12467 ( .A(n31291), .Y(n24068) );
  INVX1 U12468 ( .A(n24068), .Y(n24069) );
  BUFX2 U12469 ( .A(n31310), .Y(n24070) );
  BUFX2 U12470 ( .A(n31327), .Y(n24071) );
  BUFX2 U12471 ( .A(n31347), .Y(n24072) );
  BUFX2 U12472 ( .A(n31367), .Y(n24073) );
  BUFX2 U12473 ( .A(n31387), .Y(n24074) );
  BUFX2 U12474 ( .A(n31407), .Y(n24075) );
  BUFX2 U12475 ( .A(n31428), .Y(n24076) );
  INVX1 U12476 ( .A(n31448), .Y(n24077) );
  INVX1 U12477 ( .A(n24077), .Y(n24078) );
  BUFX2 U12478 ( .A(n31467), .Y(n24079) );
  INVX1 U12479 ( .A(n31472), .Y(n24080) );
  INVX1 U12480 ( .A(n24080), .Y(n24081) );
  INVX1 U12481 ( .A(n31487), .Y(n24082) );
  INVX1 U12482 ( .A(n24082), .Y(n24083) );
  INVX1 U12483 ( .A(n31491), .Y(n24084) );
  INVX1 U12484 ( .A(n24084), .Y(n24085) );
  INVX1 U12485 ( .A(n31510), .Y(n24086) );
  INVX1 U12486 ( .A(n24086), .Y(n24087) );
  INVX1 U12487 ( .A(n31524), .Y(n24088) );
  INVX1 U12488 ( .A(n24088), .Y(n24089) );
  INVX1 U12489 ( .A(n31529), .Y(n24090) );
  INVX1 U12490 ( .A(n24090), .Y(n24091) );
  BUFX2 U12491 ( .A(n31549), .Y(n24092) );
  INVX1 U12492 ( .A(n31569), .Y(n24093) );
  INVX1 U12493 ( .A(n24093), .Y(n24094) );
  INVX1 U12494 ( .A(n31590), .Y(n24095) );
  INVX1 U12495 ( .A(n24095), .Y(n24096) );
  INVX1 U12496 ( .A(n31609), .Y(n24097) );
  INVX1 U12497 ( .A(n24097), .Y(n24098) );
  INVX1 U12498 ( .A(n31629), .Y(n24099) );
  INVX1 U12499 ( .A(n24099), .Y(n24100) );
  INVX1 U12500 ( .A(n31645), .Y(n24101) );
  INVX1 U12501 ( .A(n24101), .Y(n24102) );
  INVX1 U12502 ( .A(n31684), .Y(n24103) );
  INVX1 U12503 ( .A(n24103), .Y(n24104) );
  BUFX2 U12504 ( .A(n31723), .Y(n24105) );
  INVX1 U12505 ( .A(n31743), .Y(n24106) );
  INVX1 U12506 ( .A(n24106), .Y(n24107) );
  BUFX2 U12507 ( .A(n31756), .Y(n24108) );
  BUFX2 U12508 ( .A(n31761), .Y(n24109) );
  BUFX2 U12509 ( .A(n31796), .Y(n24110) );
  INVX1 U12510 ( .A(n31801), .Y(n24111) );
  INVX1 U12511 ( .A(n24111), .Y(n24112) );
  BUFX2 U12512 ( .A(n31835), .Y(n24113) );
  INVX1 U12513 ( .A(n31840), .Y(n24114) );
  INVX1 U12514 ( .A(n24114), .Y(n24115) );
  INVX1 U12515 ( .A(n31860), .Y(n24116) );
  INVX1 U12516 ( .A(n24116), .Y(n24117) );
  INVX1 U12517 ( .A(n31875), .Y(n24118) );
  INVX1 U12518 ( .A(n24118), .Y(n24119) );
  INVX1 U12519 ( .A(n31881), .Y(n24120) );
  INVX1 U12520 ( .A(n24120), .Y(n24121) );
  INVX1 U12521 ( .A(n32552), .Y(n24122) );
  INVX1 U12522 ( .A(n24122), .Y(n24123) );
  INVX1 U12523 ( .A(n21145), .Y(n24124) );
  INVX1 U12524 ( .A(n32919), .Y(n24125) );
  INVX1 U12525 ( .A(n24125), .Y(n24126) );
  INVX1 U12526 ( .A(n33027), .Y(n24127) );
  BUFX2 U12527 ( .A(n33476), .Y(n24128) );
  BUFX2 U12528 ( .A(n33479), .Y(n24129) );
  BUFX2 U12529 ( .A(n33482), .Y(n24130) );
  BUFX2 U12530 ( .A(n33486), .Y(n24131) );
  BUFX2 U12531 ( .A(n33509), .Y(n24132) );
  BUFX2 U12532 ( .A(n33522), .Y(n24133) );
  BUFX2 U12533 ( .A(n33525), .Y(n24134) );
  BUFX2 U12534 ( .A(n33528), .Y(n24135) );
  BUFX2 U12535 ( .A(n33535), .Y(n24136) );
  BUFX2 U12536 ( .A(n33542), .Y(n24137) );
  BUFX2 U12537 ( .A(n33677), .Y(n24138) );
  BUFX2 U12538 ( .A(n33692), .Y(n24139) );
  BUFX2 U12539 ( .A(n33699), .Y(n24140) );
  BUFX2 U12540 ( .A(n33714), .Y(n24141) );
  BUFX2 U12541 ( .A(n33721), .Y(n24142) );
  BUFX2 U12542 ( .A(n33736), .Y(n24143) );
  BUFX2 U12543 ( .A(n33742), .Y(n24144) );
  BUFX2 U12544 ( .A(n33758), .Y(n24145) );
  BUFX2 U12545 ( .A(n33765), .Y(n24146) );
  BUFX2 U12546 ( .A(n33780), .Y(n24147) );
  BUFX2 U12547 ( .A(n33787), .Y(n24148) );
  BUFX2 U12548 ( .A(n33799), .Y(n24149) );
  BUFX2 U12549 ( .A(n33802), .Y(n24150) );
  BUFX2 U12550 ( .A(n33805), .Y(n24151) );
  BUFX2 U12551 ( .A(n33809), .Y(n24152) );
  BUFX2 U12552 ( .A(n33822), .Y(n24153) );
  BUFX2 U12553 ( .A(n33825), .Y(n24154) );
  BUFX2 U12554 ( .A(n33828), .Y(n24155) );
  BUFX2 U12555 ( .A(n33832), .Y(n24156) );
  BUFX2 U12556 ( .A(n33845), .Y(n24157) );
  BUFX2 U12557 ( .A(n33848), .Y(n24158) );
  BUFX2 U12558 ( .A(n33851), .Y(n24159) );
  BUFX2 U12559 ( .A(n33855), .Y(n24160) );
  BUFX2 U12560 ( .A(n33868), .Y(n24161) );
  BUFX2 U12561 ( .A(n33871), .Y(n24162) );
  BUFX2 U12562 ( .A(n33874), .Y(n24163) );
  BUFX2 U12563 ( .A(n33878), .Y(n24164) );
  BUFX2 U12564 ( .A(n33893), .Y(n24165) );
  BUFX2 U12565 ( .A(n33896), .Y(n24166) );
  BUFX2 U12566 ( .A(n33899), .Y(n24167) );
  BUFX2 U12567 ( .A(n33903), .Y(n24168) );
  BUFX2 U12568 ( .A(n33907), .Y(n24169) );
  INVX4 U12569 ( .A(n29354), .Y(n29360) );
  BUFX2 U12570 ( .A(n33911), .Y(n24170) );
  INVX4 U12571 ( .A(n29343), .Y(n29350) );
  BUFX2 U12572 ( .A(n29694), .Y(n24171) );
  BUFX2 U12573 ( .A(n30069), .Y(n24172) );
  BUFX2 U12574 ( .A(n30693), .Y(n24173) );
  BUFX2 U12575 ( .A(n30712), .Y(n24174) );
  BUFX2 U12576 ( .A(n30732), .Y(n24175) );
  BUFX2 U12577 ( .A(n30752), .Y(n24176) );
  BUFX2 U12578 ( .A(n30772), .Y(n24177) );
  BUFX2 U12579 ( .A(n30792), .Y(n24178) );
  BUFX2 U12580 ( .A(n30812), .Y(n24179) );
  BUFX2 U12581 ( .A(n30832), .Y(n24180) );
  BUFX2 U12582 ( .A(n30852), .Y(n24181) );
  BUFX2 U12583 ( .A(n30872), .Y(n24182) );
  BUFX2 U12584 ( .A(n30893), .Y(n24183) );
  BUFX2 U12585 ( .A(n30913), .Y(n24184) );
  BUFX2 U12586 ( .A(n30933), .Y(n24185) );
  BUFX2 U12587 ( .A(n30953), .Y(n24186) );
  BUFX2 U12588 ( .A(n30974), .Y(n24187) );
  BUFX2 U12589 ( .A(n30994), .Y(n24188) );
  BUFX2 U12590 ( .A(n31010), .Y(n24189) );
  BUFX2 U12591 ( .A(n31031), .Y(n24190) );
  BUFX2 U12592 ( .A(n31048), .Y(n24191) );
  BUFX2 U12593 ( .A(n31069), .Y(n24192) );
  BUFX2 U12594 ( .A(n31088), .Y(n24193) );
  BUFX2 U12595 ( .A(n31109), .Y(n24194) );
  BUFX2 U12596 ( .A(n31128), .Y(n24195) );
  BUFX2 U12597 ( .A(n31149), .Y(n24196) );
  BUFX2 U12598 ( .A(n31166), .Y(n24197) );
  BUFX2 U12599 ( .A(n31186), .Y(n24198) );
  BUFX2 U12600 ( .A(n31205), .Y(n24199) );
  BUFX2 U12601 ( .A(n31226), .Y(n24200) );
  BUFX2 U12602 ( .A(n31245), .Y(n24201) );
  BUFX2 U12603 ( .A(n31266), .Y(n24202) );
  BUFX2 U12604 ( .A(n31284), .Y(n24203) );
  BUFX2 U12605 ( .A(n31302), .Y(n24204) );
  BUFX2 U12606 ( .A(n31320), .Y(n24205) );
  BUFX2 U12607 ( .A(n31339), .Y(n24206) );
  BUFX2 U12608 ( .A(n31360), .Y(n24207) );
  BUFX2 U12609 ( .A(n31379), .Y(n24208) );
  BUFX2 U12610 ( .A(n31400), .Y(n24209) );
  BUFX2 U12611 ( .A(n31420), .Y(n24210) );
  BUFX2 U12612 ( .A(n31441), .Y(n24211) );
  BUFX2 U12613 ( .A(n31459), .Y(n24212) );
  BUFX2 U12614 ( .A(n31480), .Y(n24213) );
  BUFX2 U12615 ( .A(n31498), .Y(n24214) );
  BUFX2 U12616 ( .A(n31517), .Y(n24215) );
  BUFX2 U12617 ( .A(n31536), .Y(n24216) );
  BUFX2 U12618 ( .A(n31557), .Y(n24217) );
  BUFX2 U12619 ( .A(n31577), .Y(n24218) );
  BUFX2 U12620 ( .A(n31597), .Y(n24219) );
  BUFX2 U12621 ( .A(n31617), .Y(n24220) );
  BUFX2 U12622 ( .A(n31634), .Y(n24221) );
  BUFX2 U12623 ( .A(n31653), .Y(n24222) );
  BUFX2 U12624 ( .A(n31671), .Y(n24223) );
  BUFX2 U12625 ( .A(n31691), .Y(n24224) );
  BUFX2 U12626 ( .A(n31710), .Y(n24225) );
  BUFX2 U12627 ( .A(n31731), .Y(n24226) );
  BUFX2 U12628 ( .A(n31748), .Y(n24227) );
  BUFX2 U12629 ( .A(n31769), .Y(n24228) );
  BUFX2 U12630 ( .A(n31788), .Y(n24229) );
  BUFX2 U12631 ( .A(n31808), .Y(n24230) );
  BUFX2 U12632 ( .A(n31827), .Y(n24231) );
  BUFX2 U12633 ( .A(n31847), .Y(n24232) );
  BUFX2 U12634 ( .A(n31866), .Y(n24233) );
  BUFX2 U12635 ( .A(n31889), .Y(n24234) );
  BUFX2 U12636 ( .A(n32189), .Y(n24235) );
  INVX4 U12637 ( .A(n29319), .Y(n29318) );
  INVX1 U12638 ( .A(n34430), .Y(n24236) );
  INVX1 U12639 ( .A(n24236), .Y(n24237) );
  AND2X2 U12640 ( .A(n25913), .B(n32204), .Y(n30704) );
  INVX1 U12641 ( .A(n30704), .Y(n24238) );
  AND2X2 U12642 ( .A(n25917), .B(n32219), .Y(n30764) );
  INVX1 U12643 ( .A(n30764), .Y(n24239) );
  AND2X2 U12644 ( .A(n25919), .B(n32224), .Y(n30783) );
  INVX1 U12645 ( .A(n30783), .Y(n24240) );
  AND2X2 U12646 ( .A(n25920), .B(n32229), .Y(n30804) );
  INVX1 U12647 ( .A(n30804), .Y(n24241) );
  AND2X2 U12648 ( .A(n29224), .B(n26714), .Y(n30818) );
  INVX1 U12649 ( .A(n21441), .Y(n24242) );
  INVX1 U12650 ( .A(n24242), .Y(n24243) );
  INVX1 U12651 ( .A(n30103), .Y(n30443) );
  INVX1 U12652 ( .A(n25129), .Y(n31851) );
  INVX1 U12653 ( .A(n34336), .Y(n24244) );
  INVX1 U12654 ( .A(n24244), .Y(n24245) );
  BUFX2 U12655 ( .A(n29623), .Y(n24246) );
  BUFX2 U12656 ( .A(n15196), .Y(n24247) );
  AND2X2 U12657 ( .A(n26078), .B(n25404), .Y(n29876) );
  INVX1 U12658 ( .A(n29876), .Y(n24248) );
  AND2X2 U12659 ( .A(n21217), .B(net114546), .Y(n33177) );
  INVX1 U12660 ( .A(n33177), .Y(n24249) );
  AND2X2 U12661 ( .A(n23441), .B(net114546), .Y(n33179) );
  INVX1 U12662 ( .A(n33179), .Y(n24250) );
  AND2X2 U12663 ( .A(n26339), .B(net114546), .Y(n33189) );
  INVX1 U12664 ( .A(n33189), .Y(n24251) );
  AND2X2 U12665 ( .A(n21183), .B(net114546), .Y(n33192) );
  INVX1 U12666 ( .A(n33192), .Y(n24252) );
  AND2X1 U12667 ( .A(T[5]), .B(n16224), .Y(n16218) );
  INVX1 U12668 ( .A(n16218), .Y(n24253) );
  AND2X1 U12669 ( .A(T[5]), .B(n16143), .Y(n16137) );
  INVX1 U12670 ( .A(n16137), .Y(n24254) );
  AND2X1 U12671 ( .A(T[5]), .B(n15992), .Y(n15986) );
  INVX1 U12672 ( .A(n15986), .Y(n24255) );
  BUFX2 U12673 ( .A(n29556), .Y(n24256) );
  BUFX2 U12674 ( .A(n29884), .Y(n24257) );
  BUFX2 U12675 ( .A(n29899), .Y(n24258) );
  BUFX2 U12676 ( .A(n33159), .Y(n24259) );
  INVX1 U12677 ( .A(n34337), .Y(n24260) );
  INVX1 U12678 ( .A(n24260), .Y(n24261) );
  INVX1 U12679 ( .A(n24263), .Y(n24262) );
  BUFX2 U12680 ( .A(n34412), .Y(n24263) );
  INVX1 U12681 ( .A(n34439), .Y(n24264) );
  INVX1 U12682 ( .A(n24264), .Y(n24265) );
  AND2X2 U12683 ( .A(n27256), .B(n29508), .Y(n25114) );
  INVX1 U12684 ( .A(n25114), .Y(n24266) );
  AND2X1 U12685 ( .A(n16143), .B(n29661), .Y(n16136) );
  INVX1 U12686 ( .A(n16136), .Y(n24267) );
  AND2X1 U12687 ( .A(n15992), .B(n29682), .Y(n15985) );
  INVX1 U12688 ( .A(n15985), .Y(n24268) );
  AND2X2 U12689 ( .A(invdirect_s2[2]), .B(n33993), .Y(n30634) );
  INVX1 U12690 ( .A(n30634), .Y(n24269) );
  AND2X2 U12691 ( .A(invdirect_s2[1]), .B(n33993), .Y(n30654) );
  INVX1 U12692 ( .A(n30654), .Y(n24270) );
  BUFX2 U12693 ( .A(n30060), .Y(n24271) );
  INVX1 U12694 ( .A(n15566), .Y(n24272) );
  INVX1 U12695 ( .A(n24272), .Y(n24273) );
  INVX1 U12696 ( .A(n15535), .Y(n24274) );
  INVX1 U12697 ( .A(n24274), .Y(n24275) );
  INVX1 U12698 ( .A(n15222), .Y(n24276) );
  INVX1 U12699 ( .A(n24276), .Y(n24277) );
  BUFX2 U12700 ( .A(n15918), .Y(n24278) );
  INVX1 U12701 ( .A(n29748), .Y(n24279) );
  OR2X2 U12702 ( .A(n22968), .B(n25397), .Y(n30478) );
  INVX1 U12703 ( .A(n30478), .Y(n24280) );
  INVX1 U12704 ( .A(n14372), .Y(n24281) );
  INVX1 U12705 ( .A(n25328), .Y(n24282) );
  INVX1 U12706 ( .A(n29691), .Y(n24283) );
  AND2X2 U12707 ( .A(n29414), .B(n25438), .Y(n33444) );
  INVX1 U12708 ( .A(n33444), .Y(n24284) );
  AND2X2 U12709 ( .A(n29390), .B(n25438), .Y(n33449) );
  INVX1 U12710 ( .A(n33449), .Y(n24285) );
  AND2X2 U12711 ( .A(n29390), .B(n25427), .Y(n33472) );
  INVX1 U12712 ( .A(n33472), .Y(n24286) );
  AND2X2 U12713 ( .A(n29414), .B(n25426), .Y(n33489) );
  INVX1 U12714 ( .A(n33489), .Y(n24287) );
  AND2X2 U12715 ( .A(n29390), .B(n25426), .Y(n33495) );
  INVX1 U12716 ( .A(n33495), .Y(n24288) );
  AND2X2 U12717 ( .A(n29390), .B(n25457), .Y(n33518) );
  INVX1 U12718 ( .A(n33518), .Y(n24289) );
  INVX4 U12719 ( .A(n29392), .Y(n29390) );
  AND2X2 U12720 ( .A(n29390), .B(n25424), .Y(n33574) );
  INVX1 U12721 ( .A(n33574), .Y(n24290) );
  AND2X2 U12722 ( .A(n29389), .B(n25432), .Y(n33596) );
  INVX1 U12723 ( .A(n33596), .Y(n24291) );
  AND2X2 U12724 ( .A(n29389), .B(n26940), .Y(n33618) );
  INVX1 U12725 ( .A(n33618), .Y(n24292) );
  AND2X2 U12726 ( .A(n29389), .B(n25440), .Y(n33640) );
  INVX1 U12727 ( .A(n33640), .Y(n24293) );
  AND2X2 U12728 ( .A(n29389), .B(n33682), .Y(n33683) );
  INVX1 U12729 ( .A(n33683), .Y(n24294) );
  AND2X2 U12730 ( .A(n29388), .B(n26942), .Y(n33705) );
  INVX1 U12731 ( .A(n33705), .Y(n24295) );
  AND2X2 U12732 ( .A(n29388), .B(n26765), .Y(n33727) );
  INVX1 U12733 ( .A(n33727), .Y(n24296) );
  AND2X2 U12734 ( .A(n29388), .B(n23111), .Y(n33749) );
  INVX1 U12735 ( .A(n33749), .Y(n24297) );
  AND2X2 U12736 ( .A(n29388), .B(n21378), .Y(n33771) );
  INVX1 U12737 ( .A(n33771), .Y(n24298) );
  INVX4 U12738 ( .A(n29393), .Y(n29388) );
  AND2X2 U12739 ( .A(n29388), .B(n27021), .Y(n33816) );
  INVX1 U12740 ( .A(n33816), .Y(n24299) );
  AND2X2 U12741 ( .A(n29387), .B(n21375), .Y(n33838) );
  INVX1 U12742 ( .A(n33838), .Y(n24300) );
  AND2X2 U12743 ( .A(n26058), .B(n23432), .Y(n34371) );
  INVX1 U12744 ( .A(n34371), .Y(n24301) );
  BUFX2 U12745 ( .A(n30058), .Y(n24302) );
  AND2X2 U12746 ( .A(n25455), .B(n25452), .Y(n29905) );
  INVX1 U12747 ( .A(n29905), .Y(n24303) );
  AND2X2 U12748 ( .A(n25426), .B(n25351), .Y(n29915) );
  INVX1 U12749 ( .A(n29915), .Y(n24304) );
  AND2X2 U12750 ( .A(n25427), .B(n25347), .Y(n29926) );
  INVX1 U12751 ( .A(n29926), .Y(n24305) );
  AND2X2 U12752 ( .A(n25438), .B(n25350), .Y(n29936) );
  INVX1 U12753 ( .A(n29936), .Y(n24306) );
  AND2X2 U12754 ( .A(n25773), .B(n25353), .Y(n29949) );
  INVX1 U12755 ( .A(n29949), .Y(n24307) );
  AND2X2 U12756 ( .A(n21384), .B(n21435), .Y(n29959) );
  INVX1 U12757 ( .A(n29959), .Y(n24308) );
  AND2X2 U12758 ( .A(n33368), .B(n25453), .Y(n29971) );
  INVX1 U12759 ( .A(n29971), .Y(n24309) );
  AND2X2 U12760 ( .A(n33338), .B(n25355), .Y(n29982) );
  INVX1 U12761 ( .A(n29982), .Y(n24310) );
  AND2X2 U12762 ( .A(n25429), .B(n25442), .Y(n29994) );
  INVX1 U12763 ( .A(n29994), .Y(n24311) );
  AND2X2 U12764 ( .A(n25430), .B(n26269), .Y(n30005) );
  INVX1 U12765 ( .A(n30005), .Y(n24312) );
  AND2X2 U12766 ( .A(n33246), .B(n23112), .Y(n30015) );
  INVX1 U12767 ( .A(n30015), .Y(n24313) );
  AND2X2 U12768 ( .A(n21387), .B(n27195), .Y(n30028) );
  INVX1 U12769 ( .A(n30028), .Y(n24314) );
  AND2X2 U12770 ( .A(n34323), .B(n33140), .Y(n33141) );
  INVX1 U12771 ( .A(n33141), .Y(n24315) );
  AND2X2 U12772 ( .A(n21538), .B(n23602), .Y(n34202) );
  INVX1 U12773 ( .A(n34202), .Y(n24316) );
  BUFX2 U12774 ( .A(n33093), .Y(n24317) );
  BUFX2 U12775 ( .A(n33138), .Y(n24318) );
  INVX1 U12776 ( .A(n34299), .Y(n24319) );
  INVX1 U12777 ( .A(n24319), .Y(n24320) );
  BUFX2 U12778 ( .A(n34370), .Y(n24321) );
  BUFX2 U12779 ( .A(n34388), .Y(n24322) );
  BUFX2 U12780 ( .A(n16071), .Y(n24323) );
  AND2X2 U12781 ( .A(T[0]), .B(n23095), .Y(n25328) );
  INVX1 U12782 ( .A(n25328), .Y(n24324) );
  BUFX2 U12783 ( .A(n30059), .Y(n24325) );
  INVX1 U12784 ( .A(n33149), .Y(n24326) );
  INVX1 U12785 ( .A(n24326), .Y(n24327) );
  AND2X2 U12786 ( .A(n29509), .B(n29508), .Y(n29514) );
  INVX1 U12787 ( .A(n29514), .Y(n24328) );
  INVX1 U12788 ( .A(n29596), .Y(n24329) );
  INVX1 U12789 ( .A(n30692), .Y(n24330) );
  INVX1 U12790 ( .A(n24330), .Y(n24331) );
  INVX1 U12791 ( .A(n30711), .Y(n24332) );
  INVX1 U12792 ( .A(n24332), .Y(n24333) );
  BUFX2 U12793 ( .A(n30731), .Y(n24334) );
  INVX1 U12794 ( .A(n30751), .Y(n24335) );
  INVX1 U12795 ( .A(n24335), .Y(n24336) );
  INVX1 U12796 ( .A(n30771), .Y(n24337) );
  INVX1 U12797 ( .A(n24337), .Y(n24338) );
  INVX1 U12798 ( .A(n30791), .Y(n24339) );
  INVX1 U12799 ( .A(n24339), .Y(n24340) );
  INVX1 U12800 ( .A(n30811), .Y(n24341) );
  INVX1 U12801 ( .A(n24341), .Y(n24342) );
  INVX1 U12802 ( .A(n30831), .Y(n24343) );
  INVX1 U12803 ( .A(n24343), .Y(n24344) );
  INVX1 U12804 ( .A(n30851), .Y(n24345) );
  INVX1 U12805 ( .A(n24345), .Y(n24346) );
  INVX1 U12806 ( .A(n30871), .Y(n24347) );
  INVX1 U12807 ( .A(n24347), .Y(n24348) );
  INVX1 U12808 ( .A(n30892), .Y(n24349) );
  INVX1 U12809 ( .A(n24349), .Y(n24350) );
  INVX1 U12810 ( .A(n30912), .Y(n24351) );
  INVX1 U12811 ( .A(n24351), .Y(n24352) );
  INVX1 U12812 ( .A(n30932), .Y(n24353) );
  INVX1 U12813 ( .A(n24353), .Y(n24354) );
  INVX1 U12814 ( .A(n30952), .Y(n24355) );
  INVX1 U12815 ( .A(n24355), .Y(n24356) );
  INVX1 U12816 ( .A(n30973), .Y(n24357) );
  INVX1 U12817 ( .A(n24357), .Y(n24358) );
  INVX1 U12818 ( .A(n30993), .Y(n24359) );
  INVX1 U12819 ( .A(n24359), .Y(n24360) );
  INVX1 U12820 ( .A(n31009), .Y(n24361) );
  INVX1 U12821 ( .A(n24361), .Y(n24362) );
  INVX1 U12822 ( .A(n31030), .Y(n24363) );
  INVX1 U12823 ( .A(n24363), .Y(n24364) );
  INVX1 U12824 ( .A(n31047), .Y(n24365) );
  INVX1 U12825 ( .A(n24365), .Y(n24366) );
  INVX1 U12826 ( .A(n31068), .Y(n24367) );
  INVX1 U12827 ( .A(n24367), .Y(n24368) );
  INVX1 U12828 ( .A(n31087), .Y(n24369) );
  INVX1 U12829 ( .A(n24369), .Y(n24370) );
  INVX1 U12830 ( .A(n31108), .Y(n24371) );
  INVX1 U12831 ( .A(n24371), .Y(n24372) );
  INVX1 U12832 ( .A(n31127), .Y(n24373) );
  INVX1 U12833 ( .A(n24373), .Y(n24374) );
  INVX1 U12834 ( .A(n31148), .Y(n24375) );
  INVX1 U12835 ( .A(n24375), .Y(n24376) );
  INVX1 U12836 ( .A(n31165), .Y(n24377) );
  INVX1 U12837 ( .A(n24377), .Y(n24378) );
  INVX1 U12838 ( .A(n31185), .Y(n24379) );
  INVX1 U12839 ( .A(n24379), .Y(n24380) );
  INVX1 U12840 ( .A(n31204), .Y(n24381) );
  INVX1 U12841 ( .A(n24381), .Y(n24382) );
  INVX1 U12842 ( .A(n31225), .Y(n24383) );
  INVX1 U12843 ( .A(n24383), .Y(n24384) );
  BUFX2 U12844 ( .A(n31244), .Y(n24385) );
  INVX1 U12845 ( .A(n31265), .Y(n24386) );
  INVX1 U12846 ( .A(n24386), .Y(n24387) );
  BUFX2 U12847 ( .A(n31283), .Y(n24388) );
  INVX1 U12848 ( .A(n31301), .Y(n24389) );
  INVX1 U12849 ( .A(n24389), .Y(n24390) );
  INVX1 U12850 ( .A(n31319), .Y(n24391) );
  INVX1 U12851 ( .A(n24391), .Y(n24392) );
  INVX1 U12852 ( .A(n31338), .Y(n24393) );
  INVX1 U12853 ( .A(n24393), .Y(n24394) );
  INVX1 U12854 ( .A(n31359), .Y(n24395) );
  INVX1 U12855 ( .A(n24395), .Y(n24396) );
  INVX1 U12856 ( .A(n31378), .Y(n24397) );
  INVX1 U12857 ( .A(n24397), .Y(n24398) );
  INVX1 U12858 ( .A(n31399), .Y(n24399) );
  INVX1 U12859 ( .A(n24399), .Y(n24400) );
  INVX1 U12860 ( .A(n31419), .Y(n24401) );
  INVX1 U12861 ( .A(n24401), .Y(n24402) );
  INVX1 U12862 ( .A(n31440), .Y(n24403) );
  INVX1 U12863 ( .A(n24403), .Y(n24404) );
  INVX1 U12864 ( .A(n31458), .Y(n24405) );
  INVX1 U12865 ( .A(n24405), .Y(n24406) );
  INVX1 U12866 ( .A(n31479), .Y(n24407) );
  INVX1 U12867 ( .A(n24407), .Y(n24408) );
  BUFX2 U12868 ( .A(n31497), .Y(n24409) );
  INVX1 U12869 ( .A(n31516), .Y(n24410) );
  INVX1 U12870 ( .A(n24410), .Y(n24411) );
  INVX1 U12871 ( .A(n31535), .Y(n24412) );
  INVX1 U12872 ( .A(n24412), .Y(n24413) );
  BUFX2 U12873 ( .A(n31556), .Y(n24414) );
  INVX1 U12874 ( .A(n31576), .Y(n24415) );
  INVX1 U12875 ( .A(n24415), .Y(n24416) );
  INVX1 U12876 ( .A(n31596), .Y(n24417) );
  INVX1 U12877 ( .A(n24417), .Y(n24418) );
  INVX1 U12878 ( .A(n31616), .Y(n24419) );
  INVX1 U12879 ( .A(n24419), .Y(n24420) );
  BUFX2 U12880 ( .A(n31633), .Y(n24421) );
  BUFX2 U12881 ( .A(n31652), .Y(n24422) );
  BUFX2 U12882 ( .A(n31670), .Y(n24423) );
  INVX1 U12883 ( .A(n31690), .Y(n24424) );
  INVX1 U12884 ( .A(n24424), .Y(n24425) );
  BUFX2 U12885 ( .A(n31709), .Y(n24426) );
  INVX1 U12886 ( .A(n31730), .Y(n24427) );
  INVX1 U12887 ( .A(n24427), .Y(n24428) );
  BUFX2 U12888 ( .A(n31747), .Y(n24429) );
  INVX1 U12889 ( .A(n31768), .Y(n24430) );
  INVX1 U12890 ( .A(n24430), .Y(n24431) );
  BUFX2 U12891 ( .A(n31787), .Y(n24432) );
  INVX1 U12892 ( .A(n31807), .Y(n24433) );
  INVX1 U12893 ( .A(n24433), .Y(n24434) );
  BUFX2 U12894 ( .A(n31826), .Y(n24435) );
  INVX1 U12895 ( .A(n31846), .Y(n24436) );
  INVX1 U12896 ( .A(n24436), .Y(n24437) );
  BUFX2 U12897 ( .A(n31865), .Y(n24438) );
  INVX1 U12898 ( .A(n31888), .Y(n24439) );
  INVX1 U12899 ( .A(n24439), .Y(n24440) );
  BUFX2 U12900 ( .A(n29699), .Y(n24441) );
  INVX1 U12901 ( .A(n24443), .Y(n24442) );
  BUFX2 U12902 ( .A(n30048), .Y(n24443) );
  AND2X2 U12903 ( .A(n21414), .B(n29629), .Y(n29598) );
  INVX1 U12904 ( .A(n29598), .Y(n24444) );
  AND2X2 U12905 ( .A(n30038), .B(n33900), .Y(n29741) );
  INVX1 U12906 ( .A(n29741), .Y(n24445) );
  AND2X2 U12907 ( .A(n25885), .B(n25715), .Y(n30661) );
  INVX1 U12908 ( .A(n30661), .Y(n24446) );
  AND2X2 U12909 ( .A(n29224), .B(n27166), .Y(n30676) );
  AND2X2 U12910 ( .A(n25887), .B(n32199), .Y(n30681) );
  INVX1 U12911 ( .A(n30681), .Y(n24447) );
  AND2X2 U12912 ( .A(n29224), .B(n27070), .Y(n30699) );
  AND2X2 U12913 ( .A(n29224), .B(n26990), .Y(n30719) );
  AND2X2 U12914 ( .A(n25914), .B(n32209), .Y(n30724) );
  INVX1 U12915 ( .A(n30724), .Y(n24448) );
  AND2X2 U12916 ( .A(n29224), .B(n26925), .Y(n30738) );
  AND2X2 U12917 ( .A(n25916), .B(n32214), .Y(n30743) );
  INVX1 U12918 ( .A(n30743), .Y(n24449) );
  AND2X2 U12919 ( .A(n29224), .B(n26865), .Y(n30759) );
  AND2X2 U12920 ( .A(n29224), .B(n26809), .Y(n30778) );
  AND2X2 U12921 ( .A(n29224), .B(n26757), .Y(n30799) );
  AND2X2 U12922 ( .A(n29224), .B(n26681), .Y(n30839) );
  INVX1 U12923 ( .A(n30839), .Y(n24450) );
  AND2X2 U12924 ( .A(n29224), .B(n26649), .Y(n30858) );
  AND2X2 U12925 ( .A(n25911), .B(n32244), .Y(n30863) );
  INVX1 U12926 ( .A(n30863), .Y(n24451) );
  AND2X2 U12927 ( .A(n29224), .B(n26623), .Y(n30879) );
  INVX1 U12928 ( .A(n30879), .Y(n24452) );
  AND2X2 U12929 ( .A(n25884), .B(n32249), .Y(n30884) );
  INVX1 U12930 ( .A(n30884), .Y(n24453) );
  AND2X2 U12931 ( .A(n29224), .B(n27165), .Y(n30899) );
  INVX1 U12932 ( .A(n30899), .Y(n24454) );
  AND2X2 U12933 ( .A(n25881), .B(n32254), .Y(n30904) );
  INVX1 U12934 ( .A(n30904), .Y(n24455) );
  AND2X2 U12935 ( .A(n29225), .B(n27069), .Y(n30920) );
  AND2X2 U12936 ( .A(n25883), .B(n32259), .Y(n30925) );
  INVX1 U12937 ( .A(n30925), .Y(n24456) );
  AND2X2 U12938 ( .A(n29225), .B(n26924), .Y(n30939) );
  AND2X2 U12939 ( .A(n25907), .B(n32264), .Y(n30944) );
  INVX1 U12940 ( .A(n30944), .Y(n24457) );
  AND2X2 U12941 ( .A(n29225), .B(n26989), .Y(n30960) );
  INVX1 U12942 ( .A(n30960), .Y(n24458) );
  AND2X2 U12943 ( .A(n25909), .B(n32270), .Y(n30965) );
  INVX1 U12944 ( .A(n30965), .Y(n24459) );
  AND2X2 U12945 ( .A(n29225), .B(n26864), .Y(n30981) );
  INVX1 U12946 ( .A(n30981), .Y(n24460) );
  AND2X2 U12947 ( .A(n25910), .B(n32275), .Y(n30985) );
  INVX1 U12948 ( .A(n30985), .Y(n24461) );
  AND2X2 U12949 ( .A(n26030), .B(n23329), .Y(n30999) );
  INVX1 U12950 ( .A(n30999), .Y(n24462) );
  AND2X2 U12951 ( .A(n29288), .B(n27156), .Y(n31004) );
  INVX1 U12952 ( .A(n31004), .Y(n24463) );
  AND2X2 U12953 ( .A(n29225), .B(n26808), .Y(n31017) );
  AND2X2 U12954 ( .A(n25908), .B(n32283), .Y(n31022) );
  INVX1 U12955 ( .A(n31022), .Y(n24464) );
  AND2X2 U12956 ( .A(n26031), .B(n23334), .Y(n31036) );
  INVX1 U12957 ( .A(n31036), .Y(n24465) );
  AND2X2 U12958 ( .A(n29288), .B(n27057), .Y(n31042) );
  INVX1 U12959 ( .A(n31042), .Y(n24466) );
  AND2X2 U12960 ( .A(n29225), .B(n26756), .Y(n31055) );
  INVX1 U12961 ( .A(n31055), .Y(n24467) );
  AND2X2 U12962 ( .A(n25910), .B(n32291), .Y(n31060) );
  INVX1 U12963 ( .A(n31060), .Y(n24468) );
  AND2X2 U12964 ( .A(n26027), .B(n23338), .Y(n31074) );
  INVX1 U12965 ( .A(n31074), .Y(n24469) );
  AND2X2 U12966 ( .A(n29288), .B(n26977), .Y(n31081) );
  INVX1 U12967 ( .A(n31081), .Y(n24470) );
  AND2X2 U12968 ( .A(n29225), .B(n26713), .Y(n31095) );
  AND2X2 U12969 ( .A(n26032), .B(n23342), .Y(n31114) );
  INVX1 U12970 ( .A(n31114), .Y(n24471) );
  AND2X2 U12971 ( .A(n29288), .B(n26911), .Y(n31121) );
  INVX1 U12972 ( .A(n31121), .Y(n24472) );
  AND2X2 U12973 ( .A(n29225), .B(n26680), .Y(n31135) );
  INVX1 U12974 ( .A(n31135), .Y(n24473) );
  AND2X2 U12975 ( .A(n25880), .B(n32307), .Y(n31140) );
  INVX1 U12976 ( .A(n31140), .Y(n24474) );
  AND2X2 U12977 ( .A(n26031), .B(n23346), .Y(n31154) );
  INVX1 U12978 ( .A(n31154), .Y(n24475) );
  AND2X2 U12979 ( .A(n29288), .B(n27056), .Y(n31160) );
  INVX1 U12980 ( .A(n31160), .Y(n24476) );
  AND2X2 U12981 ( .A(n25879), .B(n32315), .Y(n31177) );
  INVX1 U12982 ( .A(n31177), .Y(n24477) );
  AND2X2 U12983 ( .A(n26029), .B(n23349), .Y(n31191) );
  INVX1 U12984 ( .A(n31191), .Y(n24478) );
  AND2X2 U12985 ( .A(n29288), .B(n27155), .Y(n31198) );
  INVX1 U12986 ( .A(n31198), .Y(n24479) );
  AND2X2 U12987 ( .A(n29225), .B(n26622), .Y(n31212) );
  AND2X2 U12988 ( .A(n26033), .B(n23353), .Y(n31231) );
  INVX1 U12989 ( .A(n31231), .Y(n24480) );
  AND2X2 U12990 ( .A(n29288), .B(n26910), .Y(n31238) );
  INVX1 U12991 ( .A(n31238), .Y(n24481) );
  AND2X2 U12992 ( .A(n29225), .B(n26597), .Y(n31252) );
  AND2X2 U12993 ( .A(n26030), .B(n26274), .Y(n31271) );
  INVX1 U12994 ( .A(n31271), .Y(n24482) );
  AND2X2 U12995 ( .A(n29288), .B(n26976), .Y(n31278) );
  INVX1 U12996 ( .A(n31278), .Y(n24483) );
  AND2X2 U12997 ( .A(n29223), .B(n27164), .Y(n31290) );
  INVX1 U12998 ( .A(n31290), .Y(n24484) );
  AND2X2 U12999 ( .A(n29223), .B(n27068), .Y(n31309) );
  INVX1 U13000 ( .A(n31309), .Y(n24485) );
  AND2X2 U13001 ( .A(n29223), .B(n26988), .Y(n31326) );
  INVX1 U13002 ( .A(n31326), .Y(n24486) );
  AND2X2 U13003 ( .A(n29223), .B(n26923), .Y(n31346) );
  INVX1 U13004 ( .A(n31346), .Y(n24487) );
  AND2X2 U13005 ( .A(n29223), .B(n26863), .Y(n31366) );
  INVX1 U13006 ( .A(n31366), .Y(n24488) );
  AND2X2 U13007 ( .A(n29223), .B(n26807), .Y(n31386) );
  INVX1 U13008 ( .A(n31386), .Y(n24489) );
  AND2X2 U13009 ( .A(n29223), .B(n26755), .Y(n31406) );
  INVX1 U13010 ( .A(n31406), .Y(n24490) );
  AND2X2 U13011 ( .A(n29223), .B(n26712), .Y(n31427) );
  INVX1 U13012 ( .A(n31427), .Y(n24491) );
  AND2X2 U13013 ( .A(n29223), .B(n26679), .Y(n31447) );
  INVX1 U13014 ( .A(n31447), .Y(n24492) );
  AND2X2 U13015 ( .A(n29223), .B(n26647), .Y(n31466) );
  INVX1 U13016 ( .A(n31466), .Y(n24493) );
  AND2X2 U13017 ( .A(n29223), .B(n26621), .Y(n31486) );
  INVX1 U13018 ( .A(n31486), .Y(n24494) );
  AND2X2 U13019 ( .A(n29222), .B(n27067), .Y(n31543) );
  AND2X2 U13020 ( .A(n25877), .B(n32391), .Y(n31548) );
  INVX1 U13021 ( .A(n31548), .Y(n24495) );
  AND2X2 U13022 ( .A(n29222), .B(n26987), .Y(n31563) );
  AND2X2 U13023 ( .A(n25876), .B(n32395), .Y(n31568) );
  INVX1 U13024 ( .A(n31568), .Y(n24496) );
  AND2X2 U13025 ( .A(n29222), .B(n26922), .Y(n31584) );
  AND2X2 U13026 ( .A(n25922), .B(n32399), .Y(n31589) );
  INVX1 U13027 ( .A(n31589), .Y(n24497) );
  AND2X2 U13028 ( .A(n25921), .B(n32403), .Y(n31608) );
  INVX1 U13029 ( .A(n31608), .Y(n24498) );
  AND2X2 U13030 ( .A(n26027), .B(n23394), .Y(n31622) );
  INVX1 U13031 ( .A(n31622), .Y(n24499) );
  AND2X2 U13032 ( .A(n29222), .B(n26806), .Y(n31640) );
  INVX1 U13033 ( .A(n31640), .Y(n24500) );
  AND2X2 U13034 ( .A(n25883), .B(n32411), .Y(n31644) );
  INVX1 U13035 ( .A(n31644), .Y(n24501) );
  AND2X2 U13036 ( .A(n26033), .B(n23398), .Y(n31658) );
  INVX1 U13037 ( .A(n31658), .Y(n24502) );
  AND2X2 U13038 ( .A(n29288), .B(n26909), .Y(n31665) );
  INVX1 U13039 ( .A(n31665), .Y(n24503) );
  AND2X2 U13040 ( .A(n29222), .B(n26754), .Y(n31678) );
  AND2X2 U13041 ( .A(n25918), .B(n32419), .Y(n31683) );
  INVX1 U13042 ( .A(n31683), .Y(n24504) );
  AND2X2 U13043 ( .A(n26028), .B(n23402), .Y(n31696) );
  INVX1 U13044 ( .A(n31696), .Y(n24505) );
  AND2X2 U13045 ( .A(n29288), .B(n27154), .Y(n31703) );
  INVX1 U13046 ( .A(n31703), .Y(n24506) );
  AND2X2 U13047 ( .A(n29222), .B(n26711), .Y(n31717) );
  AND2X2 U13048 ( .A(n25887), .B(n32427), .Y(n31722) );
  INVX1 U13049 ( .A(n31722), .Y(n24507) );
  AND2X2 U13050 ( .A(n26029), .B(n23406), .Y(n31736) );
  INVX1 U13051 ( .A(n31736), .Y(n24508) );
  AND2X2 U13052 ( .A(n29288), .B(n27055), .Y(n31742) );
  INVX1 U13053 ( .A(n31742), .Y(n24509) );
  AND2X2 U13054 ( .A(n29222), .B(n26678), .Y(n31755) );
  INVX1 U13055 ( .A(n31755), .Y(n24510) );
  AND2X2 U13056 ( .A(n26028), .B(n23411), .Y(n31774) );
  INVX1 U13057 ( .A(n31774), .Y(n24511) );
  AND2X2 U13058 ( .A(n29288), .B(n26908), .Y(n31781) );
  INVX1 U13059 ( .A(n31781), .Y(n24512) );
  AND2X2 U13060 ( .A(n29222), .B(n26646), .Y(n31795) );
  INVX1 U13061 ( .A(n31795), .Y(n24513) );
  AND2X2 U13062 ( .A(n25912), .B(n32442), .Y(n31800) );
  INVX1 U13063 ( .A(n31800), .Y(n24514) );
  AND2X2 U13064 ( .A(n26030), .B(n23415), .Y(n31813) );
  INVX1 U13065 ( .A(n31813), .Y(n24515) );
  AND2X2 U13066 ( .A(n29288), .B(n26974), .Y(n31820) );
  INVX1 U13067 ( .A(n31820), .Y(n24516) );
  AND2X2 U13068 ( .A(n29222), .B(n26620), .Y(n31834) );
  INVX1 U13069 ( .A(n31834), .Y(n24517) );
  AND2X2 U13070 ( .A(n25885), .B(n32450), .Y(n31839) );
  INVX1 U13071 ( .A(n31839), .Y(n24518) );
  AND2X2 U13072 ( .A(n26032), .B(n23419), .Y(n31853) );
  INVX1 U13073 ( .A(n31853), .Y(n24519) );
  AND2X2 U13074 ( .A(n29288), .B(n27054), .Y(n31859) );
  INVX1 U13075 ( .A(n31859), .Y(n24520) );
  AND2X2 U13076 ( .A(n29222), .B(n26595), .Y(n31874) );
  INVX1 U13077 ( .A(n31874), .Y(n24521) );
  AND2X2 U13078 ( .A(n25886), .B(n32457), .Y(n31880) );
  INVX1 U13079 ( .A(n31880), .Y(n24522) );
  AND2X2 U13080 ( .A(n29288), .B(n27179), .Y(n31905) );
  INVX1 U13081 ( .A(n31905), .Y(n24523) );
  AND2X2 U13082 ( .A(n29296), .B(n25357), .Y(n31919) );
  INVX1 U13083 ( .A(n31919), .Y(n24524) );
  AND2X2 U13084 ( .A(n29296), .B(n26935), .Y(n31926) );
  INVX1 U13085 ( .A(n31926), .Y(n24525) );
  AND2X2 U13086 ( .A(n29296), .B(n27090), .Y(n31931) );
  INVX1 U13087 ( .A(n31931), .Y(n24526) );
  AND2X2 U13088 ( .A(n29296), .B(n26816), .Y(n31936) );
  INVX1 U13089 ( .A(n31936), .Y(n24527) );
  AND2X2 U13090 ( .A(n29295), .B(n27088), .Y(n31941) );
  INVX1 U13091 ( .A(n31941), .Y(n24528) );
  AND2X2 U13092 ( .A(n29295), .B(n26761), .Y(n31946) );
  INVX1 U13093 ( .A(n31946), .Y(n24529) );
  AND2X2 U13094 ( .A(n29295), .B(n27002), .Y(n31951) );
  INVX1 U13095 ( .A(n31951), .Y(n24530) );
  AND2X2 U13096 ( .A(n29295), .B(n26875), .Y(n31957) );
  INVX1 U13097 ( .A(n31957), .Y(n24531) );
  AND2X2 U13098 ( .A(n29295), .B(n26716), .Y(n31962) );
  INVX1 U13099 ( .A(n31962), .Y(n24532) );
  AND2X2 U13100 ( .A(n29295), .B(n26763), .Y(n31967) );
  INVX1 U13101 ( .A(n31967), .Y(n24533) );
  AND2X2 U13102 ( .A(n29295), .B(n26937), .Y(n31972) );
  INVX1 U13103 ( .A(n31972), .Y(n24534) );
  AND2X2 U13104 ( .A(n29295), .B(n26877), .Y(n31976) );
  INVX1 U13105 ( .A(n31976), .Y(n24535) );
  AND2X2 U13106 ( .A(n29295), .B(n27004), .Y(n31981) );
  INVX1 U13107 ( .A(n31981), .Y(n24536) );
  AND2X2 U13108 ( .A(n29295), .B(n26818), .Y(n31986) );
  INVX1 U13109 ( .A(n31986), .Y(n24537) );
  AND2X2 U13110 ( .A(n29295), .B(n27094), .Y(n31992) );
  INVX1 U13111 ( .A(n31992), .Y(n24538) );
  AND2X2 U13112 ( .A(n29295), .B(n27092), .Y(n31997) );
  INVX1 U13113 ( .A(n31997), .Y(n24539) );
  AND2X2 U13114 ( .A(n29294), .B(n25358), .Y(n31999) );
  INVX1 U13115 ( .A(n31999), .Y(n24540) );
  AND2X2 U13116 ( .A(n29294), .B(n26873), .Y(n32002) );
  INVX1 U13117 ( .A(n32002), .Y(n24541) );
  AND2X2 U13118 ( .A(n29294), .B(n25359), .Y(n32004) );
  INVX1 U13119 ( .A(n32004), .Y(n24542) );
  AND2X2 U13120 ( .A(n29294), .B(n26759), .Y(n32007) );
  INVX1 U13121 ( .A(n32007), .Y(n24543) );
  AND2X2 U13122 ( .A(n29294), .B(n25360), .Y(n32010) );
  INVX1 U13123 ( .A(n32010), .Y(n24544) );
  AND2X2 U13124 ( .A(n29294), .B(n27112), .Y(n32013) );
  INVX1 U13125 ( .A(n32013), .Y(n24545) );
  AND2X2 U13126 ( .A(n29294), .B(n25361), .Y(n32016) );
  INVX1 U13127 ( .A(n32016), .Y(n24546) );
  AND2X2 U13128 ( .A(n29294), .B(n27015), .Y(n32019) );
  INVX1 U13129 ( .A(n32019), .Y(n24547) );
  AND2X2 U13130 ( .A(n29294), .B(n25362), .Y(n32022) );
  INVX1 U13131 ( .A(n32022), .Y(n24548) );
  AND2X2 U13132 ( .A(n29294), .B(n26814), .Y(n32025) );
  INVX1 U13133 ( .A(n32025), .Y(n24549) );
  AND2X2 U13134 ( .A(n29294), .B(n25342), .Y(n32028) );
  INVX1 U13135 ( .A(n32028), .Y(n24550) );
  AND2X2 U13136 ( .A(n29294), .B(n27109), .Y(n32031) );
  INVX1 U13137 ( .A(n32031), .Y(n24551) );
  AND2X2 U13138 ( .A(n29293), .B(n25363), .Y(n32034) );
  INVX1 U13139 ( .A(n32034), .Y(n24552) );
  AND2X2 U13140 ( .A(n29293), .B(n27012), .Y(n32037) );
  INVX1 U13141 ( .A(n32037), .Y(n24553) );
  AND2X2 U13142 ( .A(n29293), .B(n25364), .Y(n32040) );
  INVX1 U13143 ( .A(n32040), .Y(n24554) );
  AND2X2 U13144 ( .A(n29293), .B(n26947), .Y(n32044) );
  INVX1 U13145 ( .A(n32044), .Y(n24555) );
  AND2X2 U13146 ( .A(n29293), .B(n25365), .Y(n32048) );
  INVX1 U13147 ( .A(n32048), .Y(n24556) );
  AND2X2 U13148 ( .A(n29293), .B(n25366), .Y(n32052) );
  INVX1 U13149 ( .A(n32052), .Y(n24557) );
  AND2X2 U13150 ( .A(n29293), .B(n25367), .Y(n32056) );
  INVX1 U13151 ( .A(n32056), .Y(n24558) );
  AND2X2 U13152 ( .A(n29293), .B(n25368), .Y(n32059) );
  INVX1 U13153 ( .A(n32059), .Y(n24559) );
  AND2X2 U13154 ( .A(n29293), .B(n25369), .Y(n32063) );
  INVX1 U13155 ( .A(n32063), .Y(n24560) );
  AND2X2 U13156 ( .A(n29293), .B(n25370), .Y(n32067) );
  INVX1 U13157 ( .A(n32067), .Y(n24561) );
  AND2X2 U13158 ( .A(n29293), .B(n25371), .Y(n32071) );
  INVX1 U13159 ( .A(n32071), .Y(n24562) );
  AND2X2 U13160 ( .A(n29293), .B(n25372), .Y(n32075) );
  INVX1 U13161 ( .A(n32075), .Y(n24563) );
  AND2X2 U13162 ( .A(n29292), .B(n25373), .Y(n32079) );
  INVX1 U13163 ( .A(n32079), .Y(n24564) );
  AND2X2 U13164 ( .A(n29292), .B(n25374), .Y(n32083) );
  INVX1 U13165 ( .A(n32083), .Y(n24565) );
  AND2X2 U13166 ( .A(n29292), .B(n25375), .Y(n32087) );
  INVX1 U13167 ( .A(n32087), .Y(n24566) );
  AND2X2 U13168 ( .A(n29292), .B(n25376), .Y(n32090) );
  INVX1 U13169 ( .A(n32090), .Y(n24567) );
  AND2X2 U13170 ( .A(n29292), .B(n25377), .Y(n32094) );
  INVX1 U13171 ( .A(n32094), .Y(n24568) );
  AND2X2 U13172 ( .A(n29292), .B(n25378), .Y(n32098) );
  INVX1 U13173 ( .A(n32098), .Y(n24569) );
  AND2X2 U13174 ( .A(n29292), .B(n25379), .Y(n32104) );
  INVX1 U13175 ( .A(n32104), .Y(n24570) );
  AND2X2 U13176 ( .A(n29292), .B(n25380), .Y(n32108) );
  INVX1 U13177 ( .A(n32108), .Y(n24571) );
  AND2X2 U13178 ( .A(n29292), .B(n25381), .Y(n32111) );
  INVX1 U13179 ( .A(n32111), .Y(n24572) );
  AND2X2 U13180 ( .A(n29292), .B(n25383), .Y(n32114) );
  INVX1 U13181 ( .A(n32114), .Y(n24573) );
  AND2X2 U13182 ( .A(n29292), .B(n25384), .Y(n32117) );
  INVX1 U13183 ( .A(n32117), .Y(n24574) );
  AND2X2 U13184 ( .A(n29292), .B(n27009), .Y(n32120) );
  INVX1 U13185 ( .A(n32120), .Y(n24575) );
  AND2X2 U13186 ( .A(n29291), .B(n25385), .Y(n32123) );
  INVX1 U13187 ( .A(n32123), .Y(n24576) );
  AND2X2 U13188 ( .A(n29291), .B(n26944), .Y(n32126) );
  INVX1 U13189 ( .A(n32126), .Y(n24577) );
  AND2X2 U13190 ( .A(n29291), .B(n25386), .Y(n32129) );
  INVX1 U13191 ( .A(n32129), .Y(n24578) );
  AND2X2 U13192 ( .A(n29291), .B(n25387), .Y(n32131) );
  INVX1 U13193 ( .A(n32131), .Y(n24579) );
  AND2X2 U13194 ( .A(n29291), .B(n25388), .Y(n32134) );
  INVX1 U13195 ( .A(n32134), .Y(n24580) );
  AND2X2 U13196 ( .A(n29291), .B(n27106), .Y(n32137) );
  INVX1 U13197 ( .A(n32137), .Y(n24581) );
  AND2X2 U13198 ( .A(n29291), .B(n25389), .Y(n32140) );
  INVX1 U13199 ( .A(n32140), .Y(n24582) );
  AND2X2 U13200 ( .A(n29291), .B(n26943), .Y(n32143) );
  INVX1 U13201 ( .A(n32143), .Y(n24583) );
  AND2X2 U13202 ( .A(n29291), .B(n25390), .Y(n32146) );
  INVX1 U13203 ( .A(n32146), .Y(n24584) );
  AND2X2 U13204 ( .A(n29291), .B(n25391), .Y(n32148) );
  INVX1 U13205 ( .A(n32148), .Y(n24585) );
  AND2X2 U13206 ( .A(n29291), .B(n25392), .Y(n32151) );
  INVX1 U13207 ( .A(n32151), .Y(n24586) );
  AND2X2 U13208 ( .A(n29291), .B(n25433), .Y(n32156) );
  INVX1 U13209 ( .A(n32156), .Y(n24587) );
  AND2X2 U13210 ( .A(n23425), .B(n26145), .Y(n32188) );
  INVX1 U13211 ( .A(n32188), .Y(n24588) );
  AND2X2 U13212 ( .A(n3180), .B(n33609), .Y(n32551) );
  INVX1 U13213 ( .A(n32551), .Y(n24589) );
  INVX4 U13214 ( .A(n25431), .Y(n33609) );
  AND2X2 U13215 ( .A(n3246), .B(n32957), .Y(n32579) );
  AND2X2 U13216 ( .A(n3206), .B(n32528), .Y(n32624) );
  INVX1 U13217 ( .A(n32624), .Y(n24590) );
  AND2X2 U13218 ( .A(n32528), .B(n3211), .Y(n32816) );
  INVX1 U13219 ( .A(n32816), .Y(n24591) );
  AND2X2 U13220 ( .A(n3261), .B(n23451), .Y(n32860) );
  AND2X2 U13221 ( .A(n3247), .B(n32957), .Y(n32959) );
  AND2X2 U13222 ( .A(n3207), .B(n32528), .Y(n33015) );
  INVX1 U13223 ( .A(n33015), .Y(n24592) );
  AND2X2 U13224 ( .A(n29434), .B(n3223), .Y(n33436) );
  INVX1 U13225 ( .A(n33436), .Y(n24593) );
  AND2X2 U13226 ( .A(n29434), .B(n3221), .Y(n33439) );
  INVX1 U13227 ( .A(n33439), .Y(n24594) );
  AND2X2 U13228 ( .A(n29390), .B(n20856), .Y(n33442) );
  INVX1 U13229 ( .A(n33442), .Y(n24595) );
  AND2X2 U13230 ( .A(n29434), .B(n3217), .Y(n33454) );
  INVX1 U13231 ( .A(n33454), .Y(n24596) );
  AND2X2 U13232 ( .A(n29390), .B(n33462), .Y(n33457) );
  INVX1 U13233 ( .A(n33457), .Y(n24597) );
  AND2X2 U13234 ( .A(n29435), .B(n3215), .Y(n33460) );
  INVX1 U13235 ( .A(n33460), .Y(n24598) );
  AND2X2 U13236 ( .A(n29390), .B(n33471), .Y(n33464) );
  INVX1 U13237 ( .A(n33464), .Y(n24599) );
  AND2X2 U13238 ( .A(n29434), .B(n3211), .Y(n33477) );
  INVX1 U13239 ( .A(n33477), .Y(n24600) );
  AND2X2 U13240 ( .A(n29390), .B(n33485), .Y(n33480) );
  INVX1 U13241 ( .A(n33480), .Y(n24601) );
  AND2X2 U13242 ( .A(n29434), .B(n3209), .Y(n33483) );
  INVX1 U13243 ( .A(n33483), .Y(n24602) );
  AND2X2 U13244 ( .A(n29390), .B(n33494), .Y(n33487) );
  INVX1 U13245 ( .A(n33487), .Y(n24603) );
  AND2X2 U13246 ( .A(n29434), .B(n3205), .Y(n33500) );
  INVX1 U13247 ( .A(n33500), .Y(n24604) );
  AND2X2 U13248 ( .A(n29390), .B(n33508), .Y(n33503) );
  INVX1 U13249 ( .A(n33503), .Y(n24605) );
  AND2X2 U13250 ( .A(n29434), .B(n3203), .Y(n33506) );
  INVX1 U13251 ( .A(n33506), .Y(n24606) );
  AND2X2 U13252 ( .A(n29390), .B(n33517), .Y(n33510) );
  INVX1 U13253 ( .A(n33510), .Y(n24607) );
  AND2X2 U13254 ( .A(n29434), .B(n3199), .Y(n33523) );
  INVX1 U13255 ( .A(n33523), .Y(n24608) );
  AND2X2 U13256 ( .A(n29390), .B(n33531), .Y(n33526) );
  INVX1 U13257 ( .A(n33526), .Y(n24609) );
  AND2X2 U13258 ( .A(n29435), .B(n3197), .Y(n33529) );
  INVX1 U13259 ( .A(n33529), .Y(n24610) );
  AND2X2 U13260 ( .A(n29390), .B(n33538), .Y(n33533) );
  INVX1 U13261 ( .A(n33533), .Y(n24611) );
  AND2X2 U13262 ( .A(n29434), .B(n3195), .Y(n33536) );
  INVX1 U13263 ( .A(n33536), .Y(n24612) );
  AND2X2 U13264 ( .A(n23305), .B(n29391), .Y(n33540) );
  INVX1 U13265 ( .A(n33540), .Y(n24613) );
  AND2X2 U13266 ( .A(n29434), .B(n3193), .Y(n33543) );
  INVX1 U13267 ( .A(n33543), .Y(n24614) );
  AND2X2 U13268 ( .A(n29390), .B(n33551), .Y(n33546) );
  INVX1 U13269 ( .A(n33546), .Y(n24615) );
  AND2X2 U13270 ( .A(n29434), .B(n3191), .Y(n33549) );
  INVX1 U13271 ( .A(n33549), .Y(n24616) );
  AND2X2 U13272 ( .A(n29390), .B(n33573), .Y(n33553) );
  INVX1 U13273 ( .A(n33553), .Y(n24617) );
  AND2X2 U13274 ( .A(n29434), .B(n3187), .Y(n33579) );
  INVX1 U13275 ( .A(n33579), .Y(n24618) );
  AND2X2 U13276 ( .A(n29390), .B(n33587), .Y(n33582) );
  INVX1 U13277 ( .A(n33582), .Y(n24619) );
  AND2X2 U13278 ( .A(n29434), .B(n3185), .Y(n33585) );
  INVX1 U13279 ( .A(n33585), .Y(n24620) );
  AND2X2 U13280 ( .A(n29389), .B(n26521), .Y(n33589) );
  INVX1 U13281 ( .A(n33589), .Y(n24621) );
  AND2X2 U13282 ( .A(n29434), .B(n3181), .Y(n33601) );
  INVX1 U13283 ( .A(n33601), .Y(n24622) );
  AND2X2 U13284 ( .A(n29389), .B(n33609), .Y(n33604) );
  INVX1 U13285 ( .A(n33604), .Y(n24623) );
  AND2X2 U13286 ( .A(n29435), .B(n3179), .Y(n33607) );
  INVX1 U13287 ( .A(n33607), .Y(n24624) );
  AND2X2 U13288 ( .A(n29389), .B(n26518), .Y(n33611) );
  INVX1 U13289 ( .A(n33611), .Y(n24625) );
  AND2X2 U13290 ( .A(n29435), .B(n3175), .Y(n33623) );
  INVX1 U13291 ( .A(n33623), .Y(n24626) );
  AND2X2 U13292 ( .A(n29389), .B(n21232), .Y(n33626) );
  INVX1 U13293 ( .A(n33626), .Y(n24627) );
  AND2X2 U13294 ( .A(n29435), .B(n3173), .Y(n33629) );
  INVX1 U13295 ( .A(n33629), .Y(n24628) );
  AND2X2 U13296 ( .A(n29389), .B(n33639), .Y(n33632) );
  INVX1 U13297 ( .A(n33632), .Y(n24629) );
  AND2X2 U13298 ( .A(n29435), .B(n3169), .Y(n33645) );
  INVX1 U13299 ( .A(n33645), .Y(n24630) );
  AND2X2 U13300 ( .A(n29389), .B(n33653), .Y(n33648) );
  INVX1 U13301 ( .A(n33648), .Y(n24631) );
  AND2X2 U13302 ( .A(n29435), .B(n3167), .Y(n33651) );
  INVX1 U13303 ( .A(n33651), .Y(n24632) );
  AND2X2 U13304 ( .A(n29389), .B(n26519), .Y(n33655) );
  INVX1 U13305 ( .A(n33655), .Y(n24633) );
  AND2X2 U13306 ( .A(n29435), .B(n3163), .Y(n33667) );
  INVX1 U13307 ( .A(n33667), .Y(n24634) );
  AND2X2 U13308 ( .A(n29389), .B(n33661), .Y(n33670) );
  INVX1 U13309 ( .A(n33670), .Y(n24635) );
  AND2X2 U13310 ( .A(n29435), .B(n3161), .Y(n33673) );
  INVX1 U13311 ( .A(n33673), .Y(n24636) );
  AND2X2 U13312 ( .A(n29389), .B(n23469), .Y(n33676) );
  INVX1 U13313 ( .A(n33676), .Y(n24637) );
  AND2X2 U13314 ( .A(n29435), .B(n3157), .Y(n33688) );
  INVX1 U13315 ( .A(n33688), .Y(n24638) );
  AND2X2 U13316 ( .A(n29389), .B(n33696), .Y(n33691) );
  INVX1 U13317 ( .A(n33691), .Y(n24639) );
  AND2X2 U13318 ( .A(n29435), .B(n3155), .Y(n33694) );
  INVX1 U13319 ( .A(n33694), .Y(n24640) );
  AND2X2 U13320 ( .A(n29389), .B(n23468), .Y(n33698) );
  INVX1 U13321 ( .A(n33698), .Y(n24641) );
  AND2X2 U13322 ( .A(n29435), .B(n3151), .Y(n33710) );
  INVX1 U13323 ( .A(n33710), .Y(n24642) );
  AND2X2 U13324 ( .A(n29388), .B(n33718), .Y(n33713) );
  INVX1 U13325 ( .A(n33713), .Y(n24643) );
  AND2X2 U13326 ( .A(n29435), .B(n3149), .Y(n33716) );
  INVX1 U13327 ( .A(n33716), .Y(n24644) );
  AND2X2 U13328 ( .A(n29388), .B(n26060), .Y(n33720) );
  INVX1 U13329 ( .A(n33720), .Y(n24645) );
  AND2X2 U13330 ( .A(n29435), .B(n3145), .Y(n33732) );
  INVX1 U13331 ( .A(n33732), .Y(n24646) );
  AND2X2 U13332 ( .A(n29388), .B(n26077), .Y(n33735) );
  INVX1 U13333 ( .A(n33735), .Y(n24647) );
  AND2X2 U13334 ( .A(n29435), .B(n3143), .Y(n33738) );
  INVX1 U13335 ( .A(n33738), .Y(n24648) );
  AND2X2 U13336 ( .A(n29388), .B(n33748), .Y(n33741) );
  INVX1 U13337 ( .A(n33741), .Y(n24649) );
  AND2X2 U13338 ( .A(n29434), .B(n3139), .Y(n33754) );
  INVX1 U13339 ( .A(n33754), .Y(n24650) );
  AND2X2 U13340 ( .A(n29388), .B(n33762), .Y(n33757) );
  INVX1 U13341 ( .A(n33757), .Y(n24651) );
  AND2X2 U13342 ( .A(n29434), .B(n3137), .Y(n33760) );
  INVX1 U13343 ( .A(n33760), .Y(n24652) );
  AND2X2 U13344 ( .A(n29389), .B(n23466), .Y(n33764) );
  INVX1 U13345 ( .A(n33764), .Y(n24653) );
  AND2X2 U13346 ( .A(n29434), .B(n3133), .Y(n33776) );
  INVX1 U13347 ( .A(n33776), .Y(n24654) );
  AND2X2 U13348 ( .A(n29388), .B(n33784), .Y(n33779) );
  INVX1 U13349 ( .A(n33779), .Y(n24655) );
  AND2X2 U13350 ( .A(n29435), .B(n3131), .Y(n33782) );
  INVX1 U13351 ( .A(n33782), .Y(n24656) );
  AND2X2 U13352 ( .A(n29388), .B(n25771), .Y(n33786) );
  INVX1 U13353 ( .A(n33786), .Y(n24657) );
  AND2X2 U13354 ( .A(n29416), .B(n33806), .Y(n33798) );
  INVX1 U13355 ( .A(n33798), .Y(n24658) );
  AND2X2 U13356 ( .A(n29388), .B(n33806), .Y(n33801) );
  INVX1 U13357 ( .A(n33801), .Y(n24659) );
  AND2X2 U13358 ( .A(n29416), .B(n33815), .Y(n33804) );
  INVX1 U13359 ( .A(n33804), .Y(n24660) );
  AND2X2 U13360 ( .A(n29388), .B(n33815), .Y(n33808) );
  INVX1 U13361 ( .A(n33808), .Y(n24661) );
  AND2X2 U13362 ( .A(n29416), .B(n33829), .Y(n33821) );
  INVX1 U13363 ( .A(n33821), .Y(n24662) );
  AND2X2 U13364 ( .A(n29388), .B(n25675), .Y(n33824) );
  INVX1 U13365 ( .A(n33824), .Y(n24663) );
  AND2X2 U13366 ( .A(n29416), .B(n25830), .Y(n33827) );
  INVX1 U13367 ( .A(n33827), .Y(n24664) );
  AND2X2 U13368 ( .A(n29388), .B(n25830), .Y(n33831) );
  INVX1 U13369 ( .A(n33831), .Y(n24665) );
  AND2X2 U13370 ( .A(n29417), .B(n33852), .Y(n33844) );
  INVX1 U13371 ( .A(n33844), .Y(n24666) );
  AND2X2 U13372 ( .A(n29387), .B(n33852), .Y(n33847) );
  INVX1 U13373 ( .A(n33847), .Y(n24667) );
  AND2X2 U13374 ( .A(n29416), .B(n33861), .Y(n33850) );
  INVX1 U13375 ( .A(n33850), .Y(n24668) );
  AND2X2 U13376 ( .A(n29387), .B(n33861), .Y(n33854) );
  INVX1 U13377 ( .A(n33854), .Y(n24669) );
  AND2X2 U13378 ( .A(n29416), .B(n33875), .Y(n33867) );
  INVX1 U13379 ( .A(n33867), .Y(n24670) );
  AND2X2 U13380 ( .A(n29387), .B(n33875), .Y(n33870) );
  INVX1 U13381 ( .A(n33870), .Y(n24671) );
  AND2X2 U13382 ( .A(n29416), .B(n33884), .Y(n33873) );
  INVX1 U13383 ( .A(n33873), .Y(n24672) );
  AND2X2 U13384 ( .A(n29387), .B(n33884), .Y(n33877) );
  INVX1 U13385 ( .A(n33877), .Y(n24673) );
  AND2X2 U13386 ( .A(n29416), .B(n33900), .Y(n33892) );
  INVX1 U13387 ( .A(n33892), .Y(n24674) );
  AND2X2 U13388 ( .A(n29387), .B(n33900), .Y(n33895) );
  INVX1 U13389 ( .A(n33895), .Y(n24675) );
  AND2X2 U13390 ( .A(n29416), .B(n33908), .Y(n33898) );
  INVX1 U13391 ( .A(n33898), .Y(n24676) );
  AND2X2 U13392 ( .A(n29387), .B(n33908), .Y(n33902) );
  INVX1 U13393 ( .A(n33902), .Y(n24677) );
  AND2X2 U13394 ( .A(n27243), .B(n29417), .Y(n33906) );
  INVX1 U13395 ( .A(n33906), .Y(n24678) );
  AND2X2 U13396 ( .A(n27243), .B(n29391), .Y(n33910) );
  INVX1 U13397 ( .A(n33910), .Y(n24679) );
  AND2X2 U13398 ( .A(n29387), .B(n25774), .Y(n33914) );
  INVX1 U13399 ( .A(n33914), .Y(n24680) );
  AND2X2 U13400 ( .A(n23275), .B(n29391), .Y(n34194) );
  INVX1 U13401 ( .A(n34194), .Y(n24681) );
  AND2X2 U13402 ( .A(n23275), .B(n29417), .Y(n34207) );
  INVX1 U13403 ( .A(n34207), .Y(n24682) );
  AND2X2 U13404 ( .A(n34427), .B(n23277), .Y(n34429) );
  INVX1 U13405 ( .A(n34429), .Y(n24683) );
  BUFX2 U13406 ( .A(n29516), .Y(n24684) );
  BUFX2 U13407 ( .A(n29742), .Y(n24685) );
  INVX1 U13408 ( .A(n34175), .Y(n24686) );
  INVX1 U13409 ( .A(n24686), .Y(n24687) );
  INVX1 U13410 ( .A(n34236), .Y(n24688) );
  INVX1 U13411 ( .A(n24688), .Y(n24689) );
  INVX1 U13412 ( .A(n34368), .Y(n24690) );
  INVX1 U13413 ( .A(n24690), .Y(n24691) );
  BUFX2 U13414 ( .A(n15916), .Y(n24692) );
  OR2X1 U13415 ( .A(n15920), .B(n15921), .Y(n15919) );
  INVX1 U13416 ( .A(n15919), .Y(n24693) );
  BUFX2 U13417 ( .A(n30057), .Y(n24694) );
  AND2X2 U13418 ( .A(n2256), .B(n29510), .Y(n29512) );
  INVX1 U13419 ( .A(n29512), .Y(n24695) );
  BUFX2 U13420 ( .A(n30056), .Y(n24696) );
  BUFX2 U13421 ( .A(n29887), .Y(n24697) );
  BUFX2 U13422 ( .A(n29892), .Y(n24698) );
  BUFX2 U13423 ( .A(n29906), .Y(n24699) );
  BUFX2 U13424 ( .A(n29916), .Y(n24700) );
  BUFX2 U13425 ( .A(n29927), .Y(n24701) );
  BUFX2 U13426 ( .A(n29937), .Y(n24702) );
  BUFX2 U13427 ( .A(n29950), .Y(n24703) );
  BUFX2 U13428 ( .A(n29960), .Y(n24704) );
  BUFX2 U13429 ( .A(n29972), .Y(n24705) );
  BUFX2 U13430 ( .A(n29983), .Y(n24706) );
  BUFX2 U13431 ( .A(n29995), .Y(n24707) );
  BUFX2 U13432 ( .A(n30006), .Y(n24708) );
  BUFX2 U13433 ( .A(n30016), .Y(n24709) );
  BUFX2 U13434 ( .A(n30029), .Y(n24710) );
  INVX1 U13435 ( .A(n24712), .Y(n24711) );
  BUFX2 U13436 ( .A(n31911), .Y(n24712) );
  BUFX2 U13437 ( .A(n31918), .Y(n24713) );
  BUFX2 U13438 ( .A(n31925), .Y(n24714) );
  BUFX2 U13439 ( .A(n31930), .Y(n24715) );
  BUFX2 U13440 ( .A(n31935), .Y(n24716) );
  BUFX2 U13441 ( .A(n31940), .Y(n24717) );
  BUFX2 U13442 ( .A(n31945), .Y(n24718) );
  BUFX2 U13443 ( .A(n31950), .Y(n24719) );
  BUFX2 U13444 ( .A(n31956), .Y(n24720) );
  BUFX2 U13445 ( .A(n31961), .Y(n24721) );
  BUFX2 U13446 ( .A(n31966), .Y(n24722) );
  BUFX2 U13447 ( .A(n31971), .Y(n24723) );
  BUFX2 U13448 ( .A(n31975), .Y(n24724) );
  BUFX2 U13449 ( .A(n31980), .Y(n24725) );
  BUFX2 U13450 ( .A(n31985), .Y(n24726) );
  BUFX2 U13451 ( .A(n31991), .Y(n24727) );
  BUFX2 U13452 ( .A(n31996), .Y(n24728) );
  BUFX2 U13453 ( .A(n31998), .Y(n24729) );
  BUFX2 U13454 ( .A(n32001), .Y(n24730) );
  BUFX2 U13455 ( .A(n32003), .Y(n24731) );
  BUFX2 U13456 ( .A(n32006), .Y(n24732) );
  BUFX2 U13457 ( .A(n32009), .Y(n24733) );
  BUFX2 U13458 ( .A(n32012), .Y(n24734) );
  BUFX2 U13459 ( .A(n32015), .Y(n24735) );
  BUFX2 U13460 ( .A(n32018), .Y(n24736) );
  BUFX2 U13461 ( .A(n32021), .Y(n24737) );
  BUFX2 U13462 ( .A(n32024), .Y(n24738) );
  BUFX2 U13463 ( .A(n32027), .Y(n24739) );
  BUFX2 U13464 ( .A(n32030), .Y(n24740) );
  BUFX2 U13465 ( .A(n32033), .Y(n24741) );
  BUFX2 U13466 ( .A(n32036), .Y(n24742) );
  BUFX2 U13467 ( .A(n32039), .Y(n24743) );
  BUFX2 U13468 ( .A(n32043), .Y(n24744) );
  BUFX2 U13469 ( .A(n32047), .Y(n24745) );
  BUFX2 U13470 ( .A(n32051), .Y(n24746) );
  BUFX2 U13471 ( .A(n32055), .Y(n24747) );
  BUFX2 U13472 ( .A(n32058), .Y(n24748) );
  BUFX2 U13473 ( .A(n32062), .Y(n24749) );
  BUFX2 U13474 ( .A(n32066), .Y(n24750) );
  BUFX2 U13475 ( .A(n32070), .Y(n24751) );
  BUFX2 U13476 ( .A(n32074), .Y(n24752) );
  BUFX2 U13477 ( .A(n32078), .Y(n24753) );
  BUFX2 U13478 ( .A(n32082), .Y(n24754) );
  BUFX2 U13479 ( .A(n32086), .Y(n24755) );
  BUFX2 U13480 ( .A(n32089), .Y(n24756) );
  BUFX2 U13481 ( .A(n32093), .Y(n24757) );
  BUFX2 U13482 ( .A(n32097), .Y(n24758) );
  BUFX2 U13483 ( .A(n32103), .Y(n24759) );
  BUFX2 U13484 ( .A(n32107), .Y(n24760) );
  BUFX2 U13485 ( .A(n32110), .Y(n24761) );
  BUFX2 U13486 ( .A(n32113), .Y(n24762) );
  BUFX2 U13487 ( .A(n32116), .Y(n24763) );
  BUFX2 U13488 ( .A(n32119), .Y(n24764) );
  BUFX2 U13489 ( .A(n32122), .Y(n24765) );
  BUFX2 U13490 ( .A(n32125), .Y(n24766) );
  BUFX2 U13491 ( .A(n32128), .Y(n24767) );
  BUFX2 U13492 ( .A(n32130), .Y(n24768) );
  BUFX2 U13493 ( .A(n32133), .Y(n24769) );
  BUFX2 U13494 ( .A(n32136), .Y(n24770) );
  BUFX2 U13495 ( .A(n32139), .Y(n24771) );
  BUFX2 U13496 ( .A(n32142), .Y(n24772) );
  BUFX2 U13497 ( .A(n32145), .Y(n24773) );
  BUFX2 U13498 ( .A(n32147), .Y(n24774) );
  BUFX2 U13499 ( .A(n32150), .Y(n24775) );
  BUFX2 U13500 ( .A(n32155), .Y(n24776) );
  BUFX2 U13501 ( .A(n32187), .Y(n24777) );
  INVX1 U13502 ( .A(n32481), .Y(n24778) );
  INVX1 U13503 ( .A(n24778), .Y(n24779) );
  INVX1 U13504 ( .A(n32530), .Y(n24780) );
  INVX1 U13505 ( .A(n24780), .Y(n24781) );
  INVX1 U13506 ( .A(n32598), .Y(n24782) );
  BUFX2 U13507 ( .A(n32623), .Y(n24783) );
  INVX4 U13508 ( .A(n25452), .Y(n33517) );
  INVX1 U13509 ( .A(n32644), .Y(n24784) );
  INVX1 U13510 ( .A(n24784), .Y(n24785) );
  INVX1 U13511 ( .A(n32671), .Y(n24786) );
  INVX1 U13512 ( .A(n24786), .Y(n24787) );
  INVX1 U13513 ( .A(n32718), .Y(n24788) );
  INVX1 U13514 ( .A(n24788), .Y(n24789) );
  INVX1 U13515 ( .A(n32736), .Y(n24790) );
  INVX1 U13516 ( .A(n32815), .Y(n24791) );
  INVX1 U13517 ( .A(n24791), .Y(n24792) );
  INVX1 U13518 ( .A(n32834), .Y(n24793) );
  BUFX2 U13519 ( .A(n32905), .Y(n24794) );
  BUFX2 U13520 ( .A(n33014), .Y(n24795) );
  BUFX2 U13521 ( .A(n33435), .Y(n24796) );
  BUFX2 U13522 ( .A(n33438), .Y(n24797) );
  BUFX2 U13523 ( .A(n33441), .Y(n24798) );
  BUFX2 U13524 ( .A(n33453), .Y(n24799) );
  BUFX2 U13525 ( .A(n33456), .Y(n24800) );
  BUFX2 U13526 ( .A(n33459), .Y(n24801) );
  BUFX2 U13527 ( .A(n33463), .Y(n24802) );
  BUFX2 U13528 ( .A(n33499), .Y(n24803) );
  BUFX2 U13529 ( .A(n33502), .Y(n24804) );
  BUFX2 U13530 ( .A(n33505), .Y(n24805) );
  BUFX2 U13531 ( .A(n33532), .Y(n24806) );
  BUFX2 U13532 ( .A(n33539), .Y(n24807) );
  BUFX2 U13533 ( .A(n33545), .Y(n24808) );
  BUFX2 U13534 ( .A(n33548), .Y(n24809) );
  BUFX2 U13535 ( .A(n33552), .Y(n24810) );
  BUFX2 U13536 ( .A(n33578), .Y(n24811) );
  BUFX2 U13537 ( .A(n33581), .Y(n24812) );
  BUFX2 U13538 ( .A(n33584), .Y(n24813) );
  BUFX2 U13539 ( .A(n33588), .Y(n24814) );
  BUFX2 U13540 ( .A(n33600), .Y(n24815) );
  BUFX2 U13541 ( .A(n33603), .Y(n24816) );
  BUFX2 U13542 ( .A(n33606), .Y(n24817) );
  BUFX2 U13543 ( .A(n33610), .Y(n24818) );
  BUFX2 U13544 ( .A(n33622), .Y(n24819) );
  BUFX2 U13545 ( .A(n33625), .Y(n24820) );
  BUFX2 U13546 ( .A(n33628), .Y(n24821) );
  BUFX2 U13547 ( .A(n33631), .Y(n24822) );
  BUFX2 U13548 ( .A(n33644), .Y(n24823) );
  BUFX2 U13549 ( .A(n33647), .Y(n24824) );
  BUFX2 U13550 ( .A(n33650), .Y(n24825) );
  BUFX2 U13551 ( .A(n33654), .Y(n24826) );
  BUFX2 U13552 ( .A(n33666), .Y(n24827) );
  BUFX2 U13553 ( .A(n33669), .Y(n24828) );
  BUFX2 U13554 ( .A(n33672), .Y(n24829) );
  BUFX2 U13555 ( .A(n33687), .Y(n24830) );
  BUFX2 U13556 ( .A(n33693), .Y(n24831) );
  BUFX2 U13557 ( .A(n33709), .Y(n24832) );
  BUFX2 U13558 ( .A(n33715), .Y(n24833) );
  BUFX2 U13559 ( .A(n33731), .Y(n24834) );
  BUFX2 U13560 ( .A(n33737), .Y(n24835) );
  BUFX2 U13561 ( .A(n33753), .Y(n24836) );
  BUFX2 U13562 ( .A(n33759), .Y(n24837) );
  BUFX2 U13563 ( .A(n33775), .Y(n24838) );
  BUFX2 U13564 ( .A(n33781), .Y(n24839) );
  INVX1 U13565 ( .A(n33909), .Y(n24840) );
  INVX1 U13566 ( .A(n24840), .Y(n24841) );
  BUFX2 U13567 ( .A(n33913), .Y(n24842) );
  INVX1 U13568 ( .A(n34193), .Y(n24843) );
  INVX1 U13569 ( .A(n24843), .Y(n24844) );
  INVX1 U13570 ( .A(n34206), .Y(n24845) );
  INVX1 U13571 ( .A(n24845), .Y(n24846) );
  BUFX2 U13572 ( .A(n29877), .Y(n24847) );
  BUFX2 U13573 ( .A(n30667), .Y(n24848) );
  INVX1 U13574 ( .A(n30980), .Y(n24849) );
  INVX1 U13575 ( .A(n24849), .Y(n24850) );
  INVX1 U13576 ( .A(n31602), .Y(n24851) );
  INVX1 U13577 ( .A(n24851), .Y(n24852) );
  INVX1 U13578 ( .A(n31639), .Y(n24853) );
  INVX1 U13579 ( .A(n24853), .Y(n24854) );
  INVX1 U13580 ( .A(n34428), .Y(n24855) );
  INVX1 U13581 ( .A(n24855), .Y(n24856) );
  BUFX2 U13582 ( .A(n16214), .Y(n24857) );
  BUFX2 U13583 ( .A(n16197), .Y(n24858) );
  BUFX2 U13584 ( .A(n16133), .Y(n24859) );
  BUFX2 U13585 ( .A(n16123), .Y(n24860) );
  BUFX2 U13586 ( .A(n16116), .Y(n24861) );
  BUFX2 U13587 ( .A(n16056), .Y(n24862) );
  BUFX2 U13588 ( .A(n16039), .Y(n24863) );
  BUFX2 U13589 ( .A(n15982), .Y(n24864) );
  BUFX2 U13590 ( .A(n15972), .Y(n24865) );
  BUFX2 U13591 ( .A(n15965), .Y(n24866) );
  AND2X2 U13592 ( .A(n29624), .B(n21071), .Y(n25848) );
  INVX1 U13593 ( .A(n25848), .Y(n24867) );
  AND2X2 U13594 ( .A(n30441), .B(n29595), .Y(n29572) );
  INVX1 U13595 ( .A(n29572), .Y(n24868) );
  AND2X1 U13596 ( .A(addrLock), .B(n30064), .Y(n30065) );
  INVX1 U13597 ( .A(n30065), .Y(n24869) );
  AND2X2 U13598 ( .A(n27304), .B(n30067), .Y(n30068) );
  INVX1 U13599 ( .A(n30068), .Y(n24870) );
  INVX1 U13600 ( .A(n30077), .Y(n24871) );
  AND2X2 U13601 ( .A(n33072), .B(n23069), .Y(n33090) );
  INVX1 U13602 ( .A(n33090), .Y(n24872) );
  INVX1 U13603 ( .A(n34173), .Y(n24873) );
  OR2X2 U13604 ( .A(n34172), .B(n25346), .Y(n34173) );
  AND2X2 U13605 ( .A(n34390), .B(n25852), .Y(n34363) );
  INVX1 U13606 ( .A(n34363), .Y(n24874) );
  OR2X1 U13607 ( .A(n27192), .B(n34615), .Y(n14969) );
  INVX1 U13608 ( .A(n14969), .Y(n24875) );
  INVX1 U13609 ( .A(n14871), .Y(n24876) );
  OR2X1 U13610 ( .A(n27192), .B(n34616), .Y(n14773) );
  INVX1 U13611 ( .A(n14773), .Y(n24877) );
  BUFX2 U13612 ( .A(n29621), .Y(n24878) );
  BUFX2 U13613 ( .A(n29707), .Y(n24879) );
  INVX1 U13614 ( .A(n32776), .Y(n24882) );
  INVX1 U13615 ( .A(n24882), .Y(n24883) );
  BUFX2 U13616 ( .A(n15173), .Y(n24887) );
  INVX1 U13617 ( .A(n29753), .Y(n24888) );
  BUFX2 U13618 ( .A(n29708), .Y(n24889) );
  INVX1 U13619 ( .A(n32994), .Y(n24890) );
  INVX1 U13620 ( .A(n24890), .Y(n24891) );
  BUFX2 U13621 ( .A(n29752), .Y(n24892) );
  BUFX2 U13622 ( .A(n29763), .Y(n24893) );
  BUFX2 U13623 ( .A(n29772), .Y(n24894) );
  BUFX2 U13624 ( .A(n29780), .Y(n24895) );
  BUFX2 U13625 ( .A(n29788), .Y(n24896) );
  BUFX2 U13626 ( .A(n29797), .Y(n24897) );
  BUFX2 U13627 ( .A(n29808), .Y(n24898) );
  BUFX2 U13628 ( .A(n29818), .Y(n24899) );
  BUFX2 U13629 ( .A(n29828), .Y(n24900) );
  BUFX2 U13630 ( .A(n29839), .Y(n24901) );
  BUFX2 U13631 ( .A(n29849), .Y(n24902) );
  BUFX2 U13632 ( .A(n29857), .Y(n24903) );
  BUFX2 U13633 ( .A(n29865), .Y(n24904) );
  BUFX2 U13634 ( .A(n29874), .Y(n24905) );
  BUFX2 U13635 ( .A(n29903), .Y(n24906) );
  BUFX2 U13636 ( .A(n29913), .Y(n24907) );
  BUFX2 U13637 ( .A(n29923), .Y(n24908) );
  BUFX2 U13638 ( .A(n29934), .Y(n24909) );
  BUFX2 U13639 ( .A(n29944), .Y(n24910) );
  BUFX2 U13640 ( .A(n29957), .Y(n24911) );
  BUFX2 U13641 ( .A(n29969), .Y(n24912) );
  BUFX2 U13642 ( .A(n29980), .Y(n24913) );
  BUFX2 U13643 ( .A(n29991), .Y(n24914) );
  BUFX2 U13644 ( .A(n30003), .Y(n24915) );
  BUFX2 U13645 ( .A(n30013), .Y(n24916) );
  BUFX2 U13646 ( .A(n30025), .Y(n24917) );
  INVX1 U13647 ( .A(n32501), .Y(n24918) );
  INVX1 U13648 ( .A(n24918), .Y(n24919) );
  INVX1 U13649 ( .A(n32651), .Y(n24920) );
  INVX1 U13650 ( .A(n24920), .Y(n24921) );
  AND2X2 U13651 ( .A(n25170), .B(n25841), .Y(n14355) );
  INVX1 U13652 ( .A(n14355), .Y(n24922) );
  OR2X1 U13653 ( .A(n31868), .B(n31914), .Y(n15175) );
  INVX1 U13654 ( .A(n15175), .Y(n24923) );
  AND2X2 U13655 ( .A(n32491), .B(n23301), .Y(n27298) );
  BUFX2 U13656 ( .A(n29657), .Y(n24924) );
  AND2X2 U13657 ( .A(n2252), .B(n20813), .Y(n29473) );
  INVX1 U13658 ( .A(n29473), .Y(n24925) );
  AND2X2 U13659 ( .A(n25223), .B(n25183), .Y(n34239) );
  AND2X2 U13660 ( .A(n23200), .B(n29207), .Y(n13710) );
  INVX1 U13661 ( .A(n13710), .Y(n24926) );
  INVX1 U13662 ( .A(n13710), .Y(n24927) );
  INVX1 U13663 ( .A(n23287), .Y(n24928) );
  BUFX4 U13664 ( .A(n23110), .Y(n25332) );
  INVX1 U13665 ( .A(n23300), .Y(n24929) );
  INVX1 U13666 ( .A(n23302), .Y(n24930) );
  INVX1 U13667 ( .A(n23303), .Y(n24931) );
  BUFX2 U13668 ( .A(n14796), .Y(n24932) );
  BUFX2 U13669 ( .A(n14635), .Y(n24933) );
  BUFX2 U13670 ( .A(n14549), .Y(n24934) );
  BUFX2 U13671 ( .A(n14409), .Y(n24935) );
  AND2X2 U13672 ( .A(n25448), .B(n27254), .Y(n29660) );
  INVX1 U13673 ( .A(n29660), .Y(n24937) );
  AND2X2 U13674 ( .A(n21183), .B(n25323), .Y(n29673) );
  INVX1 U13675 ( .A(n29673), .Y(n24938) );
  AND2X2 U13676 ( .A(n29748), .B(n27252), .Y(n29724) );
  INVX1 U13677 ( .A(n29724), .Y(n24939) );
  AND2X1 U13678 ( .A(n25168), .B(n34379), .Y(n16106) );
  INVX1 U13679 ( .A(n16106), .Y(n24940) );
  AND2X2 U13680 ( .A(n29676), .B(n31917), .Y(n29680) );
  INVX1 U13681 ( .A(n29680), .Y(n24941) );
  AND2X1 U13682 ( .A(n29687), .B(n34379), .Y(n15955) );
  INVX1 U13683 ( .A(n15955), .Y(n24942) );
  INVX1 U13684 ( .A(n23304), .Y(n24943) );
  INVX1 U13685 ( .A(n23307), .Y(n24944) );
  AND2X1 U13686 ( .A(n30179), .B(n30426), .Y(n30833) );
  INVX1 U13687 ( .A(n30833), .Y(n24945) );
  AND2X1 U13688 ( .A(n30179), .B(n30440), .Y(n30873) );
  INVX1 U13689 ( .A(n30873), .Y(n24946) );
  AND2X1 U13690 ( .A(n30225), .B(n30449), .Y(n31049) );
  INVX1 U13691 ( .A(n31049), .Y(n24947) );
  AND2X1 U13692 ( .A(n30225), .B(n27311), .Y(n31089) );
  INVX1 U13693 ( .A(n31089), .Y(n24948) );
  AND2X1 U13694 ( .A(n30272), .B(n30418), .Y(n31129) );
  INVX1 U13695 ( .A(n31129), .Y(n24949) );
  AND2X1 U13696 ( .A(n30272), .B(n30432), .Y(n31167) );
  INVX1 U13697 ( .A(n31167), .Y(n24950) );
  AND2X1 U13698 ( .A(n30272), .B(n30449), .Y(n31206) );
  INVX1 U13699 ( .A(n31206), .Y(n24951) );
  AND2X1 U13700 ( .A(n30272), .B(n27311), .Y(n31246) );
  INVX1 U13701 ( .A(n31246), .Y(n24952) );
  AND2X1 U13702 ( .A(n30319), .B(n27323), .Y(n31421) );
  INVX1 U13703 ( .A(n31421), .Y(n24953) );
  AND2X1 U13704 ( .A(n27312), .B(n30426), .Y(n31460) );
  INVX1 U13705 ( .A(n31460), .Y(n24954) );
  AND2X1 U13706 ( .A(n27312), .B(n30440), .Y(n31499) );
  INVX1 U13707 ( .A(n31499), .Y(n24955) );
  AND2X1 U13708 ( .A(n30409), .B(n30449), .Y(n31672) );
  INVX1 U13709 ( .A(n31672), .Y(n24956) );
  AND2X1 U13710 ( .A(n30409), .B(n27311), .Y(n31711) );
  INVX1 U13711 ( .A(n31711), .Y(n24957) );
  AND2X1 U13712 ( .A(n30418), .B(n27324), .Y(n31749) );
  INVX1 U13713 ( .A(n31749), .Y(n24958) );
  AND2X1 U13714 ( .A(n30432), .B(n27324), .Y(n31789) );
  INVX1 U13715 ( .A(n31789), .Y(n24959) );
  AND2X1 U13716 ( .A(n30449), .B(n27324), .Y(n31828) );
  INVX1 U13717 ( .A(n31828), .Y(n24960) );
  AND2X1 U13718 ( .A(n27311), .B(n27324), .Y(n31867) );
  INVX1 U13719 ( .A(n31867), .Y(n24961) );
  INVX1 U13720 ( .A(n33157), .Y(n24962) );
  BUFX2 U13721 ( .A(n14382), .Y(n24963) );
  INVX1 U13722 ( .A(n23280), .Y(n24964) );
  AND2X1 U13723 ( .A(n27171), .B(n34351), .Y(n16139) );
  INVX1 U13724 ( .A(n16139), .Y(n24965) );
  AND2X1 U13725 ( .A(n27075), .B(n34351), .Y(n16062) );
  INVX1 U13726 ( .A(n16062), .Y(n24966) );
  AND2X2 U13727 ( .A(n29352), .B(n30499), .Y(n29774) );
  INVX1 U13728 ( .A(n29774), .Y(n24967) );
  AND2X2 U13729 ( .A(n29352), .B(n30503), .Y(n29782) );
  INVX1 U13730 ( .A(n29782), .Y(n24968) );
  AND2X2 U13731 ( .A(n29352), .B(n30518), .Y(n29810) );
  INVX1 U13732 ( .A(n29810), .Y(n24969) );
  AND2X2 U13733 ( .A(n29352), .B(n30523), .Y(n29820) );
  INVX1 U13734 ( .A(n29820), .Y(n24970) );
  AND2X2 U13735 ( .A(n29352), .B(n30527), .Y(n29830) );
  INVX1 U13736 ( .A(n29830), .Y(n24971) );
  AND2X2 U13737 ( .A(n29352), .B(n30540), .Y(n29859) );
  INVX1 U13738 ( .A(n29859), .Y(n24972) );
  INVX1 U13739 ( .A(n34174), .Y(n24973) );
  AND2X2 U13740 ( .A(n33145), .B(n33106), .Y(n33165) );
  INVX1 U13741 ( .A(n33165), .Y(n24974) );
  AND2X2 U13742 ( .A(n25424), .B(n25154), .Y(n33558) );
  INVX1 U13743 ( .A(n33558), .Y(n24975) );
  INVX1 U13744 ( .A(n23305), .Y(n24976) );
  INVX1 U13745 ( .A(n25664), .Y(n24977) );
  INVX1 U13746 ( .A(n23279), .Y(n24978) );
  AND2X2 U13747 ( .A(n25447), .B(n21007), .Y(n29665) );
  AND2X2 U13748 ( .A(n30078), .B(n29214), .Y(n30061) );
  INVX1 U13749 ( .A(n30061), .Y(n24979) );
  INVX1 U13750 ( .A(n34611), .Y(n24980) );
  INVX1 U13751 ( .A(n34611), .Y(n24981) );
  AND2X2 U13752 ( .A(n22984), .B(n23067), .Y(n34611) );
  INVX1 U13753 ( .A(n13708), .Y(n24982) );
  AND2X2 U13754 ( .A(n23280), .B(net96340), .Y(n32157) );
  INVX1 U13755 ( .A(n32157), .Y(n24983) );
  AND2X2 U13756 ( .A(n29189), .B(n34372), .Y(n25617) );
  INVX1 U13757 ( .A(n25617), .Y(n24985) );
  INVX1 U13758 ( .A(n16092), .Y(n24986) );
  INVX1 U13759 ( .A(n15941), .Y(n24987) );
  INVX1 U13760 ( .A(n21414), .Y(n29672) );
  INVX1 U13761 ( .A(n26271), .Y(n24990) );
  INVX1 U13762 ( .A(n23282), .Y(n24992) );
  INVX1 U13763 ( .A(n23285), .Y(n24993) );
  INVX1 U13764 ( .A(n23286), .Y(n24994) );
  INVX1 U13765 ( .A(n23288), .Y(n24995) );
  INVX1 U13766 ( .A(n23289), .Y(n24996) );
  INVX1 U13767 ( .A(n23291), .Y(n24997) );
  INVX1 U13768 ( .A(n23293), .Y(n24998) );
  INVX1 U13769 ( .A(n23295), .Y(n24999) );
  INVX1 U13770 ( .A(n23298), .Y(n25000) );
  INVX1 U13771 ( .A(n23299), .Y(n25001) );
  INVX1 U13772 ( .A(n23294), .Y(n25002) );
  INVX1 U13773 ( .A(n23425), .Y(n25003) );
  INVX1 U13774 ( .A(n34261), .Y(n25004) );
  INVX1 U13775 ( .A(n29590), .Y(n25005) );
  INVX1 U13776 ( .A(n23308), .Y(n25006) );
  INVX1 U13777 ( .A(n23311), .Y(n25007) );
  INVX1 U13778 ( .A(n23312), .Y(n25008) );
  INVX1 U13779 ( .A(n23313), .Y(n25009) );
  INVX1 U13780 ( .A(n23314), .Y(n25010) );
  INVX1 U13781 ( .A(n23315), .Y(n25011) );
  INVX1 U13782 ( .A(n23316), .Y(n25012) );
  INVX1 U13783 ( .A(n23317), .Y(n25013) );
  AND2X2 U13784 ( .A(n27238), .B(n30473), .Y(n31955) );
  INVX1 U13785 ( .A(n31955), .Y(n25014) );
  AND2X2 U13786 ( .A(n27246), .B(n29443), .Y(n27238) );
  INVX1 U13787 ( .A(n23318), .Y(n25015) );
  INVX1 U13788 ( .A(n23319), .Y(n25016) );
  INVX1 U13789 ( .A(n23320), .Y(n25017) );
  INVX1 U13790 ( .A(n23322), .Y(n25018) );
  INVX1 U13791 ( .A(n23323), .Y(n25019) );
  INVX1 U13792 ( .A(n23324), .Y(n25020) );
  INVX1 U13793 ( .A(n23325), .Y(n25021) );
  INVX1 U13794 ( .A(n23328), .Y(n25022) );
  INVX1 U13795 ( .A(n23330), .Y(n25023) );
  INVX1 U13796 ( .A(n23333), .Y(n25024) );
  INVX1 U13797 ( .A(n23335), .Y(n25025) );
  INVX1 U13798 ( .A(n23337), .Y(n25026) );
  INVX1 U13799 ( .A(n23339), .Y(n25027) );
  INVX1 U13800 ( .A(n23341), .Y(n25028) );
  INVX1 U13801 ( .A(n23343), .Y(n25029) );
  INVX1 U13802 ( .A(n23345), .Y(n25030) );
  INVX1 U13803 ( .A(n23348), .Y(n25031) );
  INVX1 U13804 ( .A(n23350), .Y(n25032) );
  INVX1 U13805 ( .A(n23352), .Y(n25033) );
  INVX1 U13806 ( .A(n23354), .Y(n25034) );
  INVX1 U13807 ( .A(n23356), .Y(n25035) );
  INVX1 U13808 ( .A(n23357), .Y(n25036) );
  INVX1 U13809 ( .A(n23359), .Y(n25037) );
  INVX1 U13810 ( .A(n23361), .Y(n25038) );
  INVX1 U13811 ( .A(n23363), .Y(n25039) );
  INVX1 U13812 ( .A(n23366), .Y(n25040) );
  INVX1 U13813 ( .A(n23368), .Y(n25041) );
  INVX1 U13814 ( .A(n23370), .Y(n25042) );
  INVX1 U13815 ( .A(n23372), .Y(n25043) );
  INVX1 U13816 ( .A(n23374), .Y(n25044) );
  INVX1 U13817 ( .A(n23376), .Y(n25045) );
  INVX1 U13818 ( .A(n23378), .Y(n25046) );
  INVX1 U13819 ( .A(n23380), .Y(n25047) );
  INVX1 U13820 ( .A(n23383), .Y(n25048) );
  INVX1 U13821 ( .A(n23385), .Y(n25049) );
  INVX1 U13822 ( .A(n23387), .Y(n25050) );
  INVX1 U13823 ( .A(n23389), .Y(n25051) );
  INVX1 U13824 ( .A(n23391), .Y(n25052) );
  INVX1 U13825 ( .A(n23393), .Y(n25053) );
  INVX1 U13826 ( .A(n23395), .Y(n25054) );
  INVX1 U13827 ( .A(n23397), .Y(n25055) );
  INVX1 U13828 ( .A(n23399), .Y(n25056) );
  INVX1 U13829 ( .A(n23401), .Y(n25057) );
  INVX1 U13830 ( .A(n23403), .Y(n25058) );
  INVX1 U13831 ( .A(n23405), .Y(n25059) );
  INVX1 U13832 ( .A(n23408), .Y(n25060) );
  INVX1 U13833 ( .A(n23410), .Y(n25061) );
  INVX1 U13834 ( .A(n23412), .Y(n25062) );
  INVX1 U13835 ( .A(n23414), .Y(n25063) );
  INVX1 U13836 ( .A(n23416), .Y(n25064) );
  INVX1 U13837 ( .A(n23418), .Y(n25065) );
  INVX1 U13838 ( .A(n23421), .Y(n25066) );
  INVX1 U13839 ( .A(n23423), .Y(n25067) );
  INVX1 U13840 ( .A(n23424), .Y(n25068) );
  INVX1 U13841 ( .A(n34231), .Y(n25069) );
  AND2X2 U13842 ( .A(n25706), .B(n34372), .Y(n25767) );
  INVX1 U13843 ( .A(n25767), .Y(n25070) );
  INVX1 U13844 ( .A(n25767), .Y(n25071) );
  INVX1 U13845 ( .A(n30656), .Y(n25072) );
  AND2X2 U13846 ( .A(n29352), .B(n30571), .Y(n29928) );
  INVX1 U13847 ( .A(n29928), .Y(n25073) );
  AND2X2 U13848 ( .A(n29352), .B(n30576), .Y(n29938) );
  INVX1 U13849 ( .A(n29938), .Y(n25074) );
  AND2X2 U13850 ( .A(n29352), .B(n30596), .Y(n29984) );
  INVX1 U13851 ( .A(n29984), .Y(n25075) );
  AND2X2 U13852 ( .A(n29352), .B(n30611), .Y(n30017) );
  INVX1 U13853 ( .A(n30017), .Y(n25076) );
  AND2X2 U13854 ( .A(n29352), .B(n30618), .Y(n30030) );
  INVX1 U13855 ( .A(n30030), .Y(n25077) );
  INVX1 U13856 ( .A(n21198), .Y(n25078) );
  BUFX2 U13857 ( .A(n25847), .Y(n25079) );
  INVX1 U13858 ( .A(n16281), .Y(n25080) );
  AND2X2 U13859 ( .A(n24939), .B(n27241), .Y(n29732) );
  INVX1 U13860 ( .A(n29732), .Y(n25081) );
  AND2X1 U13861 ( .A(n25623), .B(n25203), .Y(n30555) );
  INVX1 U13862 ( .A(n30555), .Y(n25082) );
  AND2X1 U13863 ( .A(n27273), .B(n29757), .Y(n30491) );
  INVX1 U13864 ( .A(n30491), .Y(n25083) );
  AND2X1 U13865 ( .A(n27273), .B(n29852), .Y(n30537) );
  INVX1 U13866 ( .A(n30537), .Y(n25084) );
  INVX1 U13867 ( .A(n23329), .Y(n25085) );
  INVX1 U13868 ( .A(n23334), .Y(n25086) );
  INVX1 U13869 ( .A(n23338), .Y(n25087) );
  INVX1 U13870 ( .A(n23342), .Y(n25088) );
  INVX1 U13871 ( .A(n23346), .Y(n25089) );
  INVX1 U13872 ( .A(n23349), .Y(n25090) );
  INVX1 U13873 ( .A(n23353), .Y(n25091) );
  INVX1 U13874 ( .A(n23394), .Y(n25092) );
  INVX1 U13875 ( .A(n23398), .Y(n25093) );
  INVX1 U13876 ( .A(n23402), .Y(n25094) );
  INVX1 U13877 ( .A(n23406), .Y(n25095) );
  INVX1 U13878 ( .A(n23411), .Y(n25096) );
  INVX1 U13879 ( .A(n23415), .Y(n25097) );
  INVX1 U13880 ( .A(n23419), .Y(n25098) );
  INVX1 U13881 ( .A(n23451), .Y(n25099) );
  INVX1 U13882 ( .A(n23281), .Y(n25100) );
  INVX1 U13883 ( .A(n32490), .Y(n25101) );
  INVX1 U13884 ( .A(n32480), .Y(n25102) );
  INVX1 U13885 ( .A(n32477), .Y(n25103) );
  INVX1 U13886 ( .A(n32478), .Y(n25104) );
  INVX1 U13887 ( .A(n23452), .Y(n25105) );
  BUFX2 U13888 ( .A(n30551), .Y(n25106) );
  AND2X1 U13889 ( .A(n30021), .B(n22942), .Y(n29746) );
  INVX1 U13890 ( .A(n29746), .Y(n25107) );
  AND2X1 U13891 ( .A(data_in[5]), .B(data_in[3]), .Y(n15174) );
  INVX1 U13892 ( .A(n15174), .Y(n25108) );
  AND2X1 U13893 ( .A(n29663), .B(n25110), .Y(n29664) );
  INVX1 U13894 ( .A(n29664), .Y(n25109) );
  INVX1 U13895 ( .A(n30441), .Y(n25110) );
  INVX1 U13896 ( .A(n29189), .Y(n25111) );
  INVX1 U13897 ( .A(n25726), .Y(n25112) );
  AND2X1 U13898 ( .A(T[1]), .B(n29667), .Y(n16117) );
  INVX1 U13899 ( .A(n16117), .Y(n25113) );
  INVX1 U13900 ( .A(n23457), .Y(n25115) );
  AND2X1 U13901 ( .A(n26837), .B(n27114), .Y(n30062) );
  INVX1 U13902 ( .A(n30062), .Y(n25116) );
  INVX1 U13903 ( .A(n29881), .Y(n25117) );
  AND2X2 U13904 ( .A(n25105), .B(n27195), .Y(n30615) );
  INVX1 U13905 ( .A(n30615), .Y(n25118) );
  OR2X2 U13906 ( .A(n34242), .B(n34250), .Y(n34248) );
  BUFX2 U13907 ( .A(n16091), .Y(n25119) );
  INVX1 U13908 ( .A(n23283), .Y(n25120) );
  INVX1 U13909 ( .A(n23284), .Y(n25121) );
  INVX1 U13910 ( .A(n23446), .Y(n25122) );
  INVX1 U13911 ( .A(n23290), .Y(n25123) );
  INVX1 U13912 ( .A(n23297), .Y(n25124) );
  INVX1 U13913 ( .A(n23449), .Y(n25125) );
  INVX1 U13914 ( .A(n25725), .Y(n25126) );
  INVX1 U13915 ( .A(n23443), .Y(n25127) );
  INVX1 U13916 ( .A(n23296), .Y(n25128) );
  AND2X2 U13917 ( .A(oc[4]), .B(n29723), .Y(n27314) );
  INVX1 U13918 ( .A(n31897), .Y(n25129) );
  BUFX2 U13919 ( .A(n33126), .Y(n25131) );
  INVX1 U13920 ( .A(n34384), .Y(n25132) );
  INVX1 U13921 ( .A(n25132), .Y(n25133) );
  AND2X2 U13922 ( .A(n25101), .B(n25452), .Y(n30561) );
  INVX1 U13923 ( .A(n30561), .Y(n25134) );
  AND2X2 U13924 ( .A(n25351), .B(n21222), .Y(n30565) );
  INVX1 U13925 ( .A(n30565), .Y(n25135) );
  AND2X2 U13926 ( .A(n25347), .B(n25155), .Y(n30570) );
  INVX1 U13927 ( .A(n30570), .Y(n25136) );
  AND2X2 U13928 ( .A(n24944), .B(n25350), .Y(n30575) );
  INVX1 U13929 ( .A(n30575), .Y(n25137) );
  AND2X2 U13930 ( .A(n25102), .B(n25353), .Y(n30580) );
  INVX1 U13931 ( .A(n30580), .Y(n25138) );
  AND2X2 U13932 ( .A(n21435), .B(n32964), .Y(n30585) );
  INVX1 U13933 ( .A(n30585), .Y(n25139) );
  AND2X2 U13934 ( .A(n25454), .B(n25444), .Y(n30590) );
  INVX1 U13935 ( .A(n30590), .Y(n25140) );
  AND2X2 U13936 ( .A(n25103), .B(n25355), .Y(n30595) );
  INVX1 U13937 ( .A(n30595), .Y(n25141) );
  AND2X2 U13938 ( .A(n25442), .B(n25394), .Y(n30600) );
  INVX1 U13939 ( .A(n30600), .Y(n25142) );
  AND2X2 U13940 ( .A(n25104), .B(n26269), .Y(n30605) );
  INVX1 U13941 ( .A(n30605), .Y(n25143) );
  AND2X2 U13942 ( .A(n25099), .B(n23112), .Y(n30610) );
  INVX1 U13943 ( .A(n30610), .Y(n25144) );
  BUFX2 U13944 ( .A(n16090), .Y(n25145) );
  BUFX2 U13945 ( .A(n15939), .Y(n25146) );
  INVX1 U13946 ( .A(n23467), .Y(n25147) );
  INVX1 U13947 ( .A(n29836), .Y(n25148) );
  INVX1 U13948 ( .A(n23450), .Y(n25149) );
  INVX1 U13949 ( .A(n33560), .Y(n25150) );
  INVX1 U13950 ( .A(n16083), .Y(n25151) );
  INVX1 U13951 ( .A(n25153), .Y(n25152) );
  BUFX2 U13952 ( .A(n29678), .Y(n25153) );
  INVX1 U13953 ( .A(n23470), .Y(n25154) );
  INVX1 U13954 ( .A(n23306), .Y(n25155) );
  AND2X1 U13955 ( .A(n25208), .B(n25422), .Y(n16084) );
  INVX1 U13956 ( .A(n16084), .Y(n25156) );
  AND2X1 U13957 ( .A(n25209), .B(n27008), .Y(n15933) );
  INVX1 U13958 ( .A(n15933), .Y(n25157) );
  INVX1 U13959 ( .A(n34256), .Y(n25158) );
  INVX1 U13960 ( .A(n25158), .Y(n25159) );
  INVX1 U13961 ( .A(n25158), .Y(n25160) );
  INVX1 U13962 ( .A(n23301), .Y(n25161) );
  INVX1 U13963 ( .A(n33158), .Y(n25162) );
  AND2X2 U13964 ( .A(n27270), .B(n30465), .Y(n31990) );
  INVX1 U13965 ( .A(n31990), .Y(n25163) );
  INVX1 U13966 ( .A(n31990), .Y(n25164) );
  AND2X2 U13967 ( .A(n27246), .B(n28220), .Y(n27270) );
  INVX1 U13968 ( .A(n23456), .Y(n25165) );
  INVX1 U13969 ( .A(n33096), .Y(n25167) );
  INVX1 U13970 ( .A(n29665), .Y(n25168) );
  INVX1 U13971 ( .A(n34317), .Y(n25169) );
  INVX1 U13972 ( .A(n30486), .Y(n25170) );
  INVX1 U13973 ( .A(net138161), .Y(net125066) );
  INVX1 U13974 ( .A(net138161), .Y(net125067) );
  INVX1 U13975 ( .A(n30910), .Y(n25171) );
  INVX1 U13976 ( .A(n30950), .Y(n25172) );
  INVX1 U13977 ( .A(n30971), .Y(n25173) );
  INVX1 U13978 ( .A(n31146), .Y(n25174) );
  INVX1 U13979 ( .A(n31183), .Y(n25175) );
  INVX1 U13980 ( .A(n31223), .Y(n25176) );
  INVX1 U13981 ( .A(n31263), .Y(n25177) );
  INVX1 U13982 ( .A(n31297), .Y(n25178) );
  INVX1 U13983 ( .A(n31357), .Y(n25179) );
  INVX1 U13984 ( .A(n31397), .Y(n25180) );
  INVX1 U13985 ( .A(n31477), .Y(n25181) );
  INVX1 U13986 ( .A(n31592), .Y(n25182) );
  INVX1 U13987 ( .A(n34243), .Y(n25183) );
  INVX1 U13988 ( .A(n30749), .Y(n25186) );
  INVX1 U13989 ( .A(n30767), .Y(n25187) );
  INVX1 U13990 ( .A(n30789), .Y(n25188) );
  INVX1 U13991 ( .A(n30829), .Y(n25189) );
  INVX1 U13992 ( .A(n31066), .Y(n25190) );
  INVX1 U13993 ( .A(n31417), .Y(n25191) );
  INVX1 U13994 ( .A(n31438), .Y(n25192) );
  INVX1 U13995 ( .A(n31766), .Y(n25193) );
  INVX1 U13996 ( .A(n25749), .Y(n25194) );
  INVX1 U13997 ( .A(n33122), .Y(n25196) );
  INVX1 U13998 ( .A(n25198), .Y(n25197) );
  BUFX2 U13999 ( .A(n16094), .Y(n25198) );
  INVX1 U14000 ( .A(n25200), .Y(n25199) );
  BUFX2 U14001 ( .A(n15943), .Y(n25200) );
  INVX1 U14002 ( .A(n34431), .Y(n25201) );
  AND2X2 U14003 ( .A(n23297), .B(n21106), .Y(n25628) );
  INVX1 U14004 ( .A(n25628), .Y(n25202) );
  INVX1 U14005 ( .A(n25628), .Y(n25203) );
  INVX1 U14006 ( .A(n33072), .Y(n25204) );
  AND2X2 U14007 ( .A(n33066), .B(n34379), .Y(n33072) );
  INVX1 U14008 ( .A(n32042), .Y(n25205) );
  INVX1 U14009 ( .A(n25855), .Y(n25206) );
  INVX1 U14010 ( .A(n16122), .Y(n25207) );
  AND2X1 U14011 ( .A(T[3]), .B(n29660), .Y(n34584) );
  INVX1 U14012 ( .A(n34584), .Y(n25208) );
  INVX1 U14013 ( .A(n34574), .Y(n25209) );
  AND2X2 U14014 ( .A(n30064), .B(n30066), .Y(n15194) );
  INVX1 U14015 ( .A(n15194), .Y(n25210) );
  INVX1 U14016 ( .A(n23309), .Y(n25211) );
  INVX1 U14017 ( .A(n23309), .Y(n25212) );
  INVX1 U14018 ( .A(n25215), .Y(n25214) );
  BUFX2 U14019 ( .A(n16212), .Y(n25215) );
  INVX1 U14020 ( .A(n16138), .Y(n25217) );
  OR2X1 U14021 ( .A(n26933), .B(n16130), .Y(n16138) );
  INVX1 U14022 ( .A(n16061), .Y(n25220) );
  OR2X1 U14023 ( .A(n27000), .B(n16053), .Y(n16061) );
  INVX1 U14024 ( .A(n34246), .Y(n25222) );
  INVX1 U14025 ( .A(n34246), .Y(n25223) );
  BUFX2 U14026 ( .A(n22998), .Y(n25224) );
  AND2X2 U14027 ( .A(n34317), .B(n23203), .Y(n34318) );
  INVX1 U14028 ( .A(n34318), .Y(n25225) );
  INVX1 U14029 ( .A(n31924), .Y(n25226) );
  INVX1 U14030 ( .A(n31924), .Y(n25227) );
  INVX1 U14031 ( .A(n31929), .Y(n25228) );
  INVX1 U14032 ( .A(n31929), .Y(n25229) );
  INVX1 U14033 ( .A(n31934), .Y(n25230) );
  INVX1 U14034 ( .A(n31934), .Y(n25231) );
  INVX1 U14035 ( .A(n31939), .Y(n25232) );
  INVX1 U14036 ( .A(n31939), .Y(n25233) );
  INVX1 U14037 ( .A(n31944), .Y(n25234) );
  INVX1 U14038 ( .A(n31944), .Y(n25235) );
  INVX1 U14039 ( .A(n31949), .Y(n25236) );
  INVX1 U14040 ( .A(n31949), .Y(n25237) );
  INVX1 U14041 ( .A(n31954), .Y(n25238) );
  INVX1 U14042 ( .A(n31954), .Y(n25239) );
  INVX1 U14043 ( .A(n31960), .Y(n25240) );
  INVX1 U14044 ( .A(n31960), .Y(n25241) );
  INVX1 U14045 ( .A(n31965), .Y(n25242) );
  INVX1 U14046 ( .A(n31965), .Y(n25243) );
  INVX1 U14047 ( .A(n31970), .Y(n25244) );
  INVX1 U14048 ( .A(n31970), .Y(n25245) );
  INVX1 U14049 ( .A(n23321), .Y(n25246) );
  INVX1 U14050 ( .A(n23321), .Y(n25247) );
  INVX1 U14051 ( .A(n31979), .Y(n25248) );
  INVX1 U14052 ( .A(n31979), .Y(n25249) );
  INVX1 U14053 ( .A(n31984), .Y(n25250) );
  INVX1 U14054 ( .A(n31984), .Y(n25251) );
  INVX1 U14055 ( .A(n31989), .Y(n25252) );
  INVX1 U14056 ( .A(n31989), .Y(n25253) );
  INVX1 U14057 ( .A(n31995), .Y(n25254) );
  INVX1 U14058 ( .A(n31995), .Y(n25255) );
  INVX1 U14059 ( .A(n23326), .Y(n25256) );
  INVX1 U14060 ( .A(n23326), .Y(n25257) );
  INVX1 U14061 ( .A(n23331), .Y(n25258) );
  INVX1 U14062 ( .A(n23331), .Y(n25259) );
  INVX1 U14063 ( .A(n32008), .Y(n25260) );
  INVX1 U14064 ( .A(n32014), .Y(n25261) );
  INVX1 U14065 ( .A(n32014), .Y(n25262) );
  INVX1 U14066 ( .A(n32020), .Y(n25263) );
  INVX1 U14067 ( .A(n32020), .Y(n25264) );
  INVX1 U14068 ( .A(n32026), .Y(n25265) );
  INVX1 U14069 ( .A(n32026), .Y(n25266) );
  INVX1 U14070 ( .A(n32032), .Y(n25267) );
  INVX1 U14071 ( .A(n32032), .Y(n25268) );
  INVX1 U14072 ( .A(n32038), .Y(n25269) );
  INVX1 U14073 ( .A(n32038), .Y(n25270) );
  INVX1 U14074 ( .A(n32046), .Y(n25271) );
  INVX1 U14075 ( .A(n32046), .Y(n25272) );
  INVX1 U14076 ( .A(n32050), .Y(n25273) );
  INVX1 U14077 ( .A(n32050), .Y(n25274) );
  INVX1 U14078 ( .A(n32054), .Y(n25275) );
  INVX1 U14079 ( .A(n32054), .Y(n25276) );
  INVX1 U14080 ( .A(n23364), .Y(n25277) );
  INVX1 U14081 ( .A(n23364), .Y(n25278) );
  INVX1 U14082 ( .A(n32061), .Y(n25279) );
  INVX1 U14083 ( .A(n32061), .Y(n25280) );
  INVX1 U14084 ( .A(n32065), .Y(n25281) );
  INVX1 U14085 ( .A(n32065), .Y(n25282) );
  INVX1 U14086 ( .A(n32069), .Y(n25283) );
  INVX1 U14087 ( .A(n32069), .Y(n25284) );
  INVX1 U14088 ( .A(n32073), .Y(n25285) );
  INVX1 U14089 ( .A(n32073), .Y(n25286) );
  INVX1 U14090 ( .A(n32077), .Y(n25287) );
  INVX1 U14091 ( .A(n32077), .Y(n25288) );
  INVX1 U14092 ( .A(n32081), .Y(n25289) );
  INVX1 U14093 ( .A(n32085), .Y(n25290) );
  INVX1 U14094 ( .A(n32085), .Y(n25291) );
  INVX1 U14095 ( .A(n23381), .Y(n25292) );
  INVX1 U14096 ( .A(n23381), .Y(n25293) );
  INVX1 U14097 ( .A(n32092), .Y(n25294) );
  INVX1 U14098 ( .A(n32092), .Y(n25295) );
  INVX1 U14099 ( .A(n32096), .Y(n25296) );
  INVX1 U14100 ( .A(n32096), .Y(n25297) );
  INVX1 U14101 ( .A(n32102), .Y(n25298) );
  INVX1 U14102 ( .A(n32102), .Y(n25299) );
  INVX1 U14103 ( .A(n32106), .Y(n25300) );
  INVX1 U14104 ( .A(n32106), .Y(n25301) );
  INVX1 U14105 ( .A(n32109), .Y(n25302) );
  INVX1 U14106 ( .A(n32109), .Y(n25303) );
  INVX1 U14107 ( .A(n32115), .Y(n25304) );
  INVX1 U14108 ( .A(n32115), .Y(n25305) );
  INVX1 U14109 ( .A(n32121), .Y(n25306) );
  INVX1 U14110 ( .A(n32121), .Y(n25307) );
  INVX1 U14111 ( .A(n32127), .Y(n25308) );
  INVX1 U14112 ( .A(n32132), .Y(n25309) );
  INVX1 U14113 ( .A(n32132), .Y(n25310) );
  INVX1 U14114 ( .A(n32138), .Y(n25311) );
  INVX1 U14115 ( .A(n32138), .Y(n25312) );
  INVX1 U14116 ( .A(n32144), .Y(n25313) );
  INVX1 U14117 ( .A(n32144), .Y(n25314) );
  INVX1 U14118 ( .A(n32149), .Y(n25315) );
  INVX1 U14119 ( .A(n32149), .Y(n25316) );
  INVX1 U14120 ( .A(n34259), .Y(n25317) );
  INVX1 U14121 ( .A(n34422), .Y(n25318) );
  INVX1 U14122 ( .A(n22988), .Y(n25319) );
  INVX1 U14123 ( .A(n34394), .Y(n25321) );
  INVX1 U14124 ( .A(n34394), .Y(n25322) );
  AND2X2 U14125 ( .A(n23645), .B(n34391), .Y(n34394) );
  AND2X2 U14126 ( .A(n29679), .B(n21183), .Y(n29670) );
  INVX1 U14127 ( .A(n29670), .Y(n25323) );
  INVX1 U14128 ( .A(n34303), .Y(n25324) );
  INVX1 U14129 ( .A(n34303), .Y(n25325) );
  INVX1 U14130 ( .A(n34241), .Y(n25326) );
  INVX1 U14131 ( .A(n34241), .Y(n25327) );
  AND2X2 U14132 ( .A(n25859), .B(T[3]), .Y(n34241) );
  BUFX2 U14133 ( .A(n33155), .Y(n25329) );
  INVX1 U14134 ( .A(n29481), .Y(n25330) );
  INVX1 U14135 ( .A(n29481), .Y(n25331) );
  INVX1 U14136 ( .A(n29583), .Y(n25333) );
  INVX1 U14137 ( .A(n25333), .Y(n25334) );
  INVX1 U14138 ( .A(n25333), .Y(n25335) );
  INVX1 U14139 ( .A(n33134), .Y(n25336) );
  INVX1 U14140 ( .A(n33134), .Y(n25337) );
  INVX1 U14141 ( .A(n21432), .Y(n25338) );
  INVX1 U14142 ( .A(n33128), .Y(n25339) );
  INVX1 U14143 ( .A(n33128), .Y(n25340) );
  AND2X1 U14144 ( .A(n29665), .B(T[0]), .Y(n34582) );
  INVX1 U14145 ( .A(n34582), .Y(n25341) );
  INVX1 U14146 ( .A(n23347), .Y(n25342) );
  INVX1 U14147 ( .A(n23428), .Y(n25344) );
  INVX1 U14148 ( .A(n23428), .Y(n25345) );
  INVX1 U14149 ( .A(n32529), .Y(n25348) );
  INVX1 U14150 ( .A(n25348), .Y(n25349) );
  INVX1 U14151 ( .A(n25348), .Y(n25350) );
  INVX1 U14152 ( .A(n32528), .Y(n25351) );
  INVX1 U14153 ( .A(n32533), .Y(n25352) );
  INVX1 U14154 ( .A(n32533), .Y(n25353) );
  INVX1 U14155 ( .A(n32536), .Y(n25354) );
  INVX1 U14156 ( .A(n32536), .Y(n25355) );
  INVX1 U14157 ( .A(n23275), .Y(n25356) );
  AND2X2 U14158 ( .A(n22941), .B(n25356), .Y(n27243) );
  AND2X2 U14159 ( .A(n22986), .B(n25356), .Y(n27241) );
  INVX1 U14160 ( .A(n23310), .Y(n25357) );
  INVX1 U14161 ( .A(n23327), .Y(n25358) );
  INVX1 U14162 ( .A(n23332), .Y(n25359) );
  INVX1 U14163 ( .A(n23336), .Y(n25360) );
  INVX1 U14164 ( .A(n23340), .Y(n25361) );
  INVX1 U14165 ( .A(n23344), .Y(n25362) );
  INVX1 U14166 ( .A(n23351), .Y(n25363) );
  INVX1 U14167 ( .A(n23355), .Y(n25364) );
  INVX1 U14168 ( .A(n23358), .Y(n25365) );
  INVX1 U14169 ( .A(n23360), .Y(n25366) );
  INVX1 U14170 ( .A(n23362), .Y(n25367) );
  INVX1 U14171 ( .A(n23365), .Y(n25368) );
  INVX1 U14172 ( .A(n23367), .Y(n25369) );
  INVX1 U14173 ( .A(n23369), .Y(n25370) );
  INVX1 U14174 ( .A(n23371), .Y(n25371) );
  INVX1 U14175 ( .A(n23373), .Y(n25372) );
  INVX1 U14176 ( .A(n23375), .Y(n25373) );
  INVX1 U14177 ( .A(n23377), .Y(n25374) );
  INVX1 U14178 ( .A(n23379), .Y(n25375) );
  INVX1 U14179 ( .A(n23382), .Y(n25376) );
  INVX1 U14180 ( .A(n23384), .Y(n25377) );
  INVX1 U14181 ( .A(n23386), .Y(n25378) );
  INVX1 U14182 ( .A(n23388), .Y(n25379) );
  INVX1 U14183 ( .A(n23390), .Y(n25380) );
  INVX1 U14184 ( .A(n23392), .Y(n25381) );
  INVX1 U14185 ( .A(n32112), .Y(n25382) );
  INVX1 U14186 ( .A(n32112), .Y(n25383) );
  INVX1 U14187 ( .A(n23396), .Y(n25384) );
  INVX1 U14188 ( .A(n23400), .Y(n25385) );
  INVX1 U14189 ( .A(n23404), .Y(n25386) );
  INVX1 U14190 ( .A(n23407), .Y(n25387) );
  INVX1 U14191 ( .A(n23409), .Y(n25388) );
  INVX1 U14192 ( .A(n23413), .Y(n25389) );
  INVX1 U14193 ( .A(n23417), .Y(n25390) );
  INVX1 U14194 ( .A(n23420), .Y(n25391) );
  INVX1 U14195 ( .A(n23422), .Y(n25392) );
  INVX1 U14196 ( .A(n32770), .Y(n25393) );
  INVX1 U14197 ( .A(n32770), .Y(n25394) );
  INVX1 U14198 ( .A(n33152), .Y(n25395) );
  INVX1 U14199 ( .A(n33152), .Y(n25396) );
  AND2X2 U14200 ( .A(n24962), .B(n25446), .Y(n33152) );
  INVX1 U14201 ( .A(n32154), .Y(n25397) );
  INVX1 U14202 ( .A(n32154), .Y(n25398) );
  INVX1 U14203 ( .A(n33167), .Y(n25399) );
  INVX1 U14204 ( .A(n25399), .Y(n25400) );
  INVX1 U14205 ( .A(n25399), .Y(n25401) );
  INVX1 U14206 ( .A(n32553), .Y(n25402) );
  INVX1 U14207 ( .A(n32553), .Y(n25403) );
  INVX1 U14208 ( .A(n32783), .Y(n25404) );
  AND2X2 U14209 ( .A(n25728), .B(T[0]), .Y(n34392) );
  INVX1 U14210 ( .A(n34392), .Y(n25405) );
  INVX1 U14211 ( .A(n29479), .Y(n25406) );
  INVX1 U14212 ( .A(n29479), .Y(n25407) );
  INVX1 U14213 ( .A(n29575), .Y(n25408) );
  INVX1 U14214 ( .A(n29575), .Y(n25409) );
  INVX1 U14215 ( .A(n31890), .Y(n25410) );
  INVX1 U14216 ( .A(n25410), .Y(n25411) );
  INVX1 U14217 ( .A(n25410), .Y(n25412) );
  INVX1 U14218 ( .A(n31899), .Y(n25413) );
  INVX1 U14219 ( .A(n25413), .Y(n25414) );
  INVX1 U14220 ( .A(n34403), .Y(n25415) );
  INVX1 U14221 ( .A(n25415), .Y(n25416) );
  INVX1 U14222 ( .A(n25415), .Y(n25417) );
  INVX1 U14223 ( .A(n33132), .Y(n25418) );
  INVX1 U14224 ( .A(n33132), .Y(n25419) );
  INVX1 U14225 ( .A(n29594), .Y(n25420) );
  AND2X2 U14226 ( .A(n27301), .B(n21007), .Y(n29594) );
  INVX1 U14227 ( .A(n29594), .Y(n25421) );
  INVX1 U14228 ( .A(n16104), .Y(n25422) );
  INVX1 U14229 ( .A(n33572), .Y(n25423) );
  INVX1 U14230 ( .A(n33572), .Y(n25424) );
  INVX1 U14231 ( .A(n33493), .Y(n25425) );
  INVX1 U14232 ( .A(n33493), .Y(n25426) );
  INVX1 U14233 ( .A(n33307), .Y(n25428) );
  INVX1 U14234 ( .A(n33307), .Y(n25429) );
  INVX1 U14235 ( .A(n33595), .Y(n25431) );
  INVX1 U14236 ( .A(n33595), .Y(n25432) );
  INVX1 U14237 ( .A(n32152), .Y(n25433) );
  INVX1 U14238 ( .A(n32152), .Y(n25434) );
  AND2X2 U14239 ( .A(n30476), .B(n30475), .Y(n32152) );
  INVX1 U14240 ( .A(n34324), .Y(n25435) );
  INVX1 U14241 ( .A(n34324), .Y(n25436) );
  INVX1 U14242 ( .A(n33448), .Y(n25437) );
  INVX1 U14243 ( .A(n33448), .Y(n25438) );
  INVX1 U14244 ( .A(n33638), .Y(n25439) );
  INVX1 U14245 ( .A(n33638), .Y(n25440) );
  INVX1 U14246 ( .A(n33002), .Y(n25442) );
  INVX1 U14247 ( .A(n32863), .Y(n25443) );
  INVX1 U14248 ( .A(n32863), .Y(n25444) );
  INVX1 U14249 ( .A(n32863), .Y(n25445) );
  AND2X2 U14250 ( .A(n29968), .B(n29331), .Y(n32863) );
  INVX1 U14251 ( .A(n32153), .Y(n25447) );
  INVX1 U14252 ( .A(n32153), .Y(n25448) );
  INVX1 U14253 ( .A(n32153), .Y(n25449) );
  AND2X2 U14254 ( .A(n29670), .B(n30410), .Y(n32153) );
  INVX1 U14255 ( .A(n8054), .Y(n25450) );
  INVX1 U14256 ( .A(n8054), .Y(n25451) );
  AND2X2 U14257 ( .A(n23477), .B(n29498), .Y(n8054) );
  AND2X2 U14258 ( .A(n23449), .B(n21106), .Y(n32910) );
  INVX1 U14259 ( .A(n32913), .Y(n25453) );
  AND2X2 U14260 ( .A(n23288), .B(n32491), .Y(n32913) );
  INVX1 U14261 ( .A(net89759), .Y(net124029) );
  INVX1 U14262 ( .A(net89759), .Y(net124030) );
  INVX1 U14263 ( .A(n33516), .Y(n25455) );
  INVX1 U14264 ( .A(n33516), .Y(n25456) );
  INVX1 U14265 ( .A(n33516), .Y(n25457) );
  AND2X2 U14266 ( .A(n23298), .B(n30626), .Y(n33516) );
  AND2X2 U14267 ( .A(n25458), .B(n25459), .Y(n21858) );
  INVX1 U14268 ( .A(n25754), .Y(n25459) );
  INVX1 U14269 ( .A(n23116), .Y(n25460) );
  NAND3X1 U14270 ( .A(n25463), .B(n25462), .C(n21177), .Y(n25464) );
  INVX1 U14271 ( .A(n33032), .Y(n25463) );
  INVX1 U14272 ( .A(n25464), .Y(n33045) );
  INVX1 U14273 ( .A(net149764), .Y(net109512) );
  MUX2X1 U14274 ( .B(n28218), .A(n28219), .S(net151429), .Y(n28217) );
  NAND3X1 U14275 ( .A(data_in[4]), .B(data_in[0]), .C(n22794), .Y(n25640) );
  INVX1 U14276 ( .A(n21162), .Y(n29384) );
  BUFX2 U14277 ( .A(grid[278]), .Y(n25465) );
  AND2X2 U14278 ( .A(n25346), .B(n29212), .Y(n25467) );
  INVX1 U14279 ( .A(n29261), .Y(n25468) );
  INVX1 U14280 ( .A(net151814), .Y(net117301) );
  AND2X2 U14281 ( .A(n9133), .B(n29378), .Y(n21790) );
  AND2X2 U14282 ( .A(n9126), .B(n29381), .Y(n21783) );
  INVX1 U14283 ( .A(n29735), .Y(n25473) );
  AND2X2 U14284 ( .A(n29269), .B(n26877), .Y(n25474) );
  INVX1 U14285 ( .A(n27105), .Y(n25475) );
  BUFX2 U14286 ( .A(grid[66]), .Y(n25478) );
  INVX1 U14287 ( .A(net112181), .Y(net117217) );
  INVX1 U14288 ( .A(n25510), .Y(n25480) );
  BUFX2 U14289 ( .A(grid[211]), .Y(n25481) );
  INVX1 U14290 ( .A(net116777), .Y(net117076) );
  NAND3X1 U14291 ( .A(n25753), .B(n27255), .C(n25647), .Y(n25483) );
  BUFX2 U14292 ( .A(grid[26]), .Y(n25484) );
  MUX2X1 U14293 ( .B(grid[358]), .A(grid[352]), .S(net149922), .Y(n28165) );
  INVX1 U14294 ( .A(n34349), .Y(n25485) );
  MUX2X1 U14295 ( .B(n28034), .A(n28033), .S(net116949), .Y(n28032) );
  BUFX2 U14296 ( .A(grid[355]), .Y(n25486) );
  BUFX2 U14297 ( .A(grid[241]), .Y(n25487) );
  BUFX2 U14298 ( .A(grid[349]), .Y(n25488) );
  INVX1 U14299 ( .A(n29627), .Y(n25489) );
  INVX1 U14300 ( .A(n13802), .Y(n29627) );
  BUFX2 U14301 ( .A(grid[253]), .Y(n25490) );
  AND2X2 U14302 ( .A(n23284), .B(n29330), .Y(n25491) );
  INVX2 U14303 ( .A(n25491), .Y(n32964) );
  BUFX2 U14304 ( .A(grid[343]), .Y(n25492) );
  BUFX2 U14305 ( .A(grid[307]), .Y(n25493) );
  BUFX2 U14306 ( .A(grid[247]), .Y(n25494) );
  BUFX2 U14307 ( .A(grid[98]), .Y(n25495) );
  BUFX2 U14308 ( .A(grid[187]), .Y(n25496) );
  BUFX2 U14309 ( .A(grid[55]), .Y(n25497) );
  BUFX2 U14310 ( .A(n25486), .Y(n25498) );
  INVX8 U14311 ( .A(net109766), .Y(net103671) );
  BUFX2 U14312 ( .A(grid[200]), .Y(n25499) );
  BUFX2 U14313 ( .A(grid[338]), .Y(n25500) );
  MUX2X1 U14314 ( .B(n27975), .A(n27960), .S(net104479), .Y(alt14_net6005) );
  MUX2X1 U14315 ( .B(n28096), .A(n28095), .S(net105822), .Y(n28094) );
  BUFX2 U14316 ( .A(grid[91]), .Y(n25501) );
  BUFX2 U14317 ( .A(grid[326]), .Y(n25502) );
  BUFX2 U14318 ( .A(grid[74]), .Y(n25503) );
  INVX1 U14319 ( .A(grid[194]), .Y(n25504) );
  INVX1 U14320 ( .A(n25504), .Y(n25505) );
  INVX1 U14321 ( .A(alt14_net96264), .Y(net116776) );
  BUFX2 U14322 ( .A(grid[265]), .Y(n25506) );
  BUFX2 U14323 ( .A(grid[43]), .Y(n25507) );
  BUFX2 U14324 ( .A(grid[38]), .Y(n25508) );
  BUFX2 U14325 ( .A(grid[230]), .Y(n25509) );
  INVX1 U14326 ( .A(net151662), .Y(net116754) );
  INVX1 U14327 ( .A(grid[37]), .Y(n25510) );
  INVX1 U14328 ( .A(n25510), .Y(n25511) );
  BUFX2 U14329 ( .A(n25497), .Y(n25512) );
  BUFX2 U14330 ( .A(grid[277]), .Y(n25513) );
  BUFX2 U14331 ( .A(n25499), .Y(n25514) );
  AND2X2 U14332 ( .A(n25466), .B(n31305), .Y(n25515) );
  BUFX2 U14333 ( .A(grid[103]), .Y(n25516) );
  MUX2X1 U14334 ( .B(grid[68]), .A(grid[62]), .S(net150133), .Y(n28090) );
  MUX2X1 U14335 ( .B(grid[248]), .A(grid[242]), .S(net137490), .Y(n28059) );
  AND2X2 U14336 ( .A(n29268), .B(n26814), .Y(n25518) );
  OR2X2 U14337 ( .A(n23456), .B(n29261), .Y(n25519) );
  NAND3X1 U14338 ( .A(n33048), .B(n33046), .C(n33047), .Y(n25528) );
  OAI21X1 U14339 ( .A(net150331), .B(net149842), .C(n30631), .Y(n25529) );
  INVX1 U14340 ( .A(n31900), .Y(n25530) );
  INVX1 U14341 ( .A(n31900), .Y(n25531) );
  INVX1 U14342 ( .A(n31900), .Y(n25532) );
  INVX1 U14343 ( .A(n31900), .Y(n25533) );
  INVX1 U14344 ( .A(n25530), .Y(n25534) );
  INVX1 U14345 ( .A(n25530), .Y(n25535) );
  INVX1 U14346 ( .A(n25530), .Y(n25536) );
  INVX1 U14347 ( .A(n25530), .Y(n25537) );
  INVX1 U14348 ( .A(n25531), .Y(n25538) );
  INVX1 U14349 ( .A(n25531), .Y(n25539) );
  INVX1 U14350 ( .A(n25531), .Y(n25540) );
  INVX1 U14351 ( .A(n25532), .Y(n25541) );
  INVX1 U14352 ( .A(n25532), .Y(n25542) );
  INVX1 U14353 ( .A(n25532), .Y(n25543) );
  INVX1 U14354 ( .A(n25532), .Y(n25544) );
  INVX1 U14355 ( .A(n25533), .Y(n25545) );
  INVX1 U14356 ( .A(n25533), .Y(n25546) );
  INVX1 U14357 ( .A(n25533), .Y(n25547) );
  BUFX2 U14358 ( .A(n25529), .Y(n25548) );
  INVX1 U14359 ( .A(n25557), .Y(n25549) );
  INVX1 U14360 ( .A(n25548), .Y(n25550) );
  INVX1 U14361 ( .A(n25548), .Y(n25551) );
  INVX1 U14362 ( .A(n25548), .Y(n25552) );
  INVX1 U14363 ( .A(n25548), .Y(n25553) );
  INVX1 U14364 ( .A(n25548), .Y(n25554) );
  INVX1 U14365 ( .A(n25556), .Y(n25555) );
  BUFX2 U14366 ( .A(n25529), .Y(n25556) );
  BUFX2 U14367 ( .A(n25529), .Y(n25557) );
  INVX1 U14368 ( .A(n25556), .Y(n25558) );
  INVX1 U14369 ( .A(n25556), .Y(n25559) );
  INVX1 U14370 ( .A(n25556), .Y(n25560) );
  INVX1 U14371 ( .A(n25556), .Y(n25561) );
  INVX1 U14372 ( .A(n25557), .Y(n25562) );
  INVX1 U14373 ( .A(n25556), .Y(n25563) );
  INVX1 U14374 ( .A(n25557), .Y(n25564) );
  INVX1 U14375 ( .A(n25557), .Y(n25565) );
  INVX1 U14376 ( .A(n25557), .Y(n25566) );
  INVX1 U14377 ( .A(n25557), .Y(n25567) );
  INVX1 U14378 ( .A(n25556), .Y(n25568) );
  INVX4 U14379 ( .A(n29264), .Y(n29261) );
  AND2X2 U14380 ( .A(n23579), .B(n21550), .Y(n27281) );
  INVX1 U14381 ( .A(n25529), .Y(n31900) );
  INVX4 U14382 ( .A(n25634), .Y(n29331) );
  INVX1 U14383 ( .A(n34187), .Y(n25569) );
  INVX1 U14384 ( .A(n27173), .Y(n25570) );
  MUX2X1 U14385 ( .B(grid[151]), .A(grid[145]), .S(net116777), .Y(n28012) );
  OR2X1 U14386 ( .A(n32803), .B(n26269), .Y(n25572) );
  INVX2 U14387 ( .A(n22677), .Y(n34317) );
  OR2X2 U14388 ( .A(n22118), .B(n32806), .Y(n32814) );
  BUFX2 U14389 ( .A(oc[28]), .Y(n25573) );
  INVX1 U14390 ( .A(n27906), .Y(n27904) );
  BUFX2 U14391 ( .A(grid[146]), .Y(n25574) );
  INVX1 U14392 ( .A(n33058), .Y(n25575) );
  BUFX2 U14393 ( .A(grid[2]), .Y(n25576) );
  BUFX2 U14394 ( .A(n25507), .Y(n25577) );
  BUFX2 U14395 ( .A(grid[73]), .Y(n25578) );
  INVX1 U14396 ( .A(n22880), .Y(n29486) );
  INVX1 U14397 ( .A(n23088), .Y(n25579) );
  INVX1 U14398 ( .A(n33175), .Y(n25580) );
  MUX2X1 U14399 ( .B(grid[31]), .A(grid[25]), .S(n26446), .Y(n28336) );
  MUX2X1 U14400 ( .B(grid[178]), .A(grid[172]), .S(n26446), .Y(n28501) );
  BUFX2 U14401 ( .A(grid[56]), .Y(n25581) );
  BUFX2 U14402 ( .A(grid[20]), .Y(n25582) );
  MUX2X1 U14403 ( .B(grid[212]), .A(grid[206]), .S(net150133), .Y(n28066) );
  MUX2X1 U14404 ( .B(grid[130]), .A(grid[124]), .S(n26446), .Y(n28507) );
  BUFX2 U14405 ( .A(n25513), .Y(n25583) );
  AND2X2 U14406 ( .A(n27272), .B(n20849), .Y(n27239) );
  MUX2X1 U14407 ( .B(grid[163]), .A(grid[157]), .S(net150220), .Y(n28013) );
  INVX2 U14408 ( .A(n26445), .Y(n26087) );
  XOR2X1 U14409 ( .A(n21112), .B(n34323), .Y(n25584) );
  XOR2X1 U14410 ( .A(n25719), .B(n25584), .Y(n34263) );
  INVX1 U14411 ( .A(net53785), .Y(net115635) );
  INVX1 U14412 ( .A(net115635), .Y(net115636) );
  BUFX2 U14413 ( .A(n34292), .Y(n25585) );
  INVX1 U14414 ( .A(net145105), .Y(net64168) );
  AND2X2 U14415 ( .A(n21544), .B(n21555), .Y(n32884) );
  INVX4 U14416 ( .A(net105778), .Y(net114151) );
  INVX1 U14417 ( .A(locTrig[2]), .Y(n25589) );
  INVX2 U14418 ( .A(n25661), .Y(n29422) );
  INVX4 U14419 ( .A(n27902), .Y(n27909) );
  MUX2X1 U14420 ( .B(grid[106]), .A(grid[100]), .S(n26517), .Y(n28510) );
  MUX2X1 U14421 ( .B(n28326), .A(n28341), .S(n33995), .Y(n28344) );
  INVX1 U14422 ( .A(n27261), .Y(n25590) );
  INVX1 U14423 ( .A(n20849), .Y(n25592) );
  AND2X2 U14424 ( .A(net149983), .B(net105822), .Y(n27244) );
  INVX2 U14425 ( .A(alt14_net96328), .Y(net105819) );
  BUFX2 U14426 ( .A(n25772), .Y(n25593) );
  INVX1 U14427 ( .A(grid[158]), .Y(n25594) );
  INVX1 U14428 ( .A(n25594), .Y(n25595) );
  AND2X2 U14429 ( .A(n29376), .B(n31169), .Y(n25596) );
  INVX1 U14430 ( .A(n33573), .Y(n25597) );
  BUFX2 U14431 ( .A(grid[266]), .Y(n25598) );
  INVX4 U14432 ( .A(net105778), .Y(net105779) );
  BUFX2 U14433 ( .A(grid[194]), .Y(n25599) );
  BUFX2 U14434 ( .A(grid[205]), .Y(n25600) );
  BUFX2 U14435 ( .A(grid[110]), .Y(n25601) );
  BUFX2 U14436 ( .A(grid[260]), .Y(n25602) );
  BUFX2 U14437 ( .A(grid[31]), .Y(n25603) );
  NOR3X1 U14438 ( .A(n23274), .B(n25111), .C(n33062), .Y(n25604) );
  INVX2 U14439 ( .A(n34369), .Y(n34395) );
  BUFX2 U14440 ( .A(grid[302]), .Y(n25605) );
  AND2X2 U14441 ( .A(n9130), .B(n21166), .Y(n21787) );
  MUX2X1 U14442 ( .B(n28054), .A(n28053), .S(net114916), .Y(n28052) );
  BUFX2 U14443 ( .A(grid[49]), .Y(n25607) );
  BUFX2 U14444 ( .A(n25511), .Y(n25608) );
  MUX2X1 U14445 ( .B(grid[322]), .A(grid[316]), .S(n21090), .Y(n28477) );
  MUX2X1 U14446 ( .B(grid[11]), .A(grid[5]), .S(n21163), .Y(n28587) );
  MUX2X1 U14447 ( .B(n28493), .A(n28492), .S(n26514), .Y(n28491) );
  MUX2X1 U14448 ( .B(grid[10]), .A(grid[4]), .S(n21097), .Y(n28525) );
  INVX1 U14449 ( .A(n13804), .Y(n34171) );
  BUFX2 U14450 ( .A(n14357), .Y(net114808) );
  INVX1 U14451 ( .A(grid[290]), .Y(n25609) );
  INVX1 U14452 ( .A(n25609), .Y(n25610) );
  INVX1 U14453 ( .A(n25620), .Y(n25611) );
  AND2X2 U14454 ( .A(n9135), .B(n29379), .Y(n21792) );
  INVX1 U14455 ( .A(n29542), .Y(n25612) );
  INVX1 U14456 ( .A(n29550), .Y(n25613) );
  INVX4 U14457 ( .A(n25439), .Y(n33653) );
  AND2X2 U14458 ( .A(n22983), .B(n22995), .Y(n25614) );
  INVX1 U14459 ( .A(n25614), .Y(n34211) );
  XNOR2X1 U14460 ( .A(n26063), .B(n34442), .Y(n34292) );
  OAI21X1 U14461 ( .A(n25863), .B(n25133), .C(n34383), .Y(n25616) );
  BUFX2 U14462 ( .A(grid[300]), .Y(n25618) );
  MUX2X1 U14463 ( .B(n28175), .A(n28178), .S(n20936), .Y(n28189) );
  MUX2X1 U14464 ( .B(n28029), .A(n28032), .S(net114244), .Y(n28036) );
  INVX1 U14465 ( .A(net150245), .Y(net114244) );
  BUFX2 U14466 ( .A(grid[61]), .Y(n25622) );
  INVX1 U14467 ( .A(n32973), .Y(n25623) );
  AND2X2 U14468 ( .A(n33053), .B(n33054), .Y(n25624) );
  AND2X2 U14469 ( .A(n30078), .B(n29215), .Y(net114546) );
  BUFX2 U14470 ( .A(grid[162]), .Y(n25625) );
  BUFX2 U14471 ( .A(grid[348]), .Y(n25626) );
  INVX1 U14472 ( .A(pLoc[3]), .Y(net114252) );
  BUFX2 U14473 ( .A(grid[276]), .Y(n25627) );
  MUX2X1 U14474 ( .B(n27993), .A(n27996), .S(net114244), .Y(n28007) );
  INVX1 U14475 ( .A(n26046), .Y(n25629) );
  INVX1 U14476 ( .A(n25629), .Y(n25630) );
  BUFX2 U14477 ( .A(grid[192]), .Y(n25631) );
  BUFX2 U14478 ( .A(grid[48]), .Y(n25632) );
  BUFX2 U14479 ( .A(grid[12]), .Y(n25633) );
  MUX2X1 U14480 ( .B(grid[82]), .A(grid[76]), .S(net105778), .Y(n28206) );
  MUX2X1 U14481 ( .B(n28201), .A(n28200), .S(net105821), .Y(n28199) );
  AND2X2 U14482 ( .A(n22996), .B(n25473), .Y(n25634) );
  BUFX2 U14483 ( .A(grid[204]), .Y(n25635) );
  BUFX2 U14484 ( .A(grid[240]), .Y(n25637) );
  INVX1 U14485 ( .A(grid[60]), .Y(n25638) );
  INVX1 U14486 ( .A(n25638), .Y(n25639) );
  AND2X2 U14487 ( .A(n30626), .B(n23288), .Y(n33617) );
  MUX2X1 U14488 ( .B(n28180), .A(n28179), .S(net105821), .Y(n28178) );
  MUX2X1 U14489 ( .B(grid[334]), .A(grid[328]), .S(net151801), .Y(n28168) );
  AND2X2 U14490 ( .A(n30626), .B(n23289), .Y(n25641) );
  INVX1 U14491 ( .A(n25641), .Y(n33338) );
  INVX1 U14492 ( .A(n21105), .Y(n25642) );
  BUFX2 U14493 ( .A(grid[252]), .Y(n25643) );
  OAI21X1 U14494 ( .A(n34322), .B(n34309), .C(n34308), .Y(n25644) );
  OR2X2 U14495 ( .A(n32947), .B(n32946), .Y(n32956) );
  INVX1 U14496 ( .A(oc[22]), .Y(n25645) );
  INVX1 U14497 ( .A(n25645), .Y(n25646) );
  INVX1 U14498 ( .A(n32704), .Y(n26070) );
  AND2X2 U14499 ( .A(n27303), .B(n29331), .Y(n27250) );
  AND2X2 U14500 ( .A(n20971), .B(n33049), .Y(n25647) );
  NAND3X1 U14501 ( .A(n25649), .B(n25604), .C(n21233), .Y(n25648) );
  INVX1 U14502 ( .A(n22997), .Y(n34362) );
  INVX4 U14503 ( .A(n34215), .Y(n29443) );
  INVX1 U14504 ( .A(n28221), .Y(n25732) );
  NOR3X1 U14505 ( .A(net110320), .B(net149850), .C(n29600), .Y(n25651) );
  INVX1 U14506 ( .A(n25651), .Y(n29697) );
  INVX1 U14507 ( .A(n30989), .Y(n25652) );
  INVX1 U14508 ( .A(net53785), .Y(net113686) );
  INVX1 U14509 ( .A(net90071), .Y(net53785) );
  BUFX2 U14510 ( .A(grid[206]), .Y(n25654) );
  BUFX2 U14511 ( .A(grid[50]), .Y(n25655) );
  BUFX2 U14512 ( .A(grid[14]), .Y(n25656) );
  INVX2 U14513 ( .A(net105821), .Y(net113308) );
  AND2X2 U14514 ( .A(n9136), .B(n29379), .Y(n21793) );
  AND2X2 U14515 ( .A(n30626), .B(n23286), .Y(n25657) );
  INVX1 U14516 ( .A(n25657), .Y(n33368) );
  AND2X2 U14517 ( .A(n30626), .B(n23296), .Y(n25658) );
  INVX1 U14518 ( .A(n25658), .Y(n33246) );
  BUFX2 U14519 ( .A(grid[62]), .Y(n25659) );
  BUFX2 U14520 ( .A(grid[242]), .Y(n25660) );
  AND2X2 U14521 ( .A(n33057), .B(n33058), .Y(n25661) );
  AND2X2 U14522 ( .A(oc[4]), .B(oc[3]), .Y(n27315) );
  INVX1 U14523 ( .A(n21028), .Y(n29491) );
  INVX2 U14524 ( .A(n20849), .Y(n26084) );
  INVX1 U14525 ( .A(n25665), .Y(n28594) );
  MUX2X1 U14526 ( .B(n28216), .A(n28215), .S(net113687), .Y(n28214) );
  INVX1 U14527 ( .A(n25690), .Y(n33125) );
  OR2X2 U14528 ( .A(n32709), .B(n32710), .Y(n32717) );
  AND2X2 U14529 ( .A(net109585), .B(n29191), .Y(n27309) );
  AND2X2 U14530 ( .A(n27304), .B(net109585), .Y(n27267) );
  INVX4 U14531 ( .A(n25437), .Y(n33462) );
  MUX2X1 U14532 ( .B(n28260), .A(n28259), .S(n26514), .Y(n28258) );
  INVX1 U14533 ( .A(net114808), .Y(net112858) );
  INVX1 U14534 ( .A(net112858), .Y(net112859) );
  MUX2X1 U14535 ( .B(n28067), .A(n28052), .S(net104479), .Y(alt14_net6130) );
  BUFX2 U14536 ( .A(n8050), .Y(n25665) );
  MUX2X1 U14537 ( .B(grid[143]), .A(grid[137]), .S(n21163), .Y(n28570) );
  MUX2X1 U14538 ( .B(grid[179]), .A(grid[173]), .S(n21097), .Y(n28563) );
  INVX1 U14539 ( .A(n34395), .Y(n25666) );
  INVX1 U14540 ( .A(n25666), .Y(n25667) );
  INVX1 U14541 ( .A(n34295), .Y(n25668) );
  OR2X2 U14542 ( .A(n8039), .B(n8038), .Y(n30045) );
  INVX1 U14543 ( .A(n31612), .Y(n25670) );
  MUX2X1 U14544 ( .B(n28051), .A(n28050), .S(net149876), .Y(n28049) );
  MUX2X1 U14545 ( .B(n28481), .A(n28480), .S(n26514), .Y(n28479) );
  INVX1 U14546 ( .A(n30639), .Y(n25672) );
  NOR3X1 U14547 ( .A(n29191), .B(n25673), .C(n25672), .Y(n25671) );
  INVX1 U14548 ( .A(n25671), .Y(n31912) );
  AND2X2 U14549 ( .A(n27304), .B(net151710), .Y(n25673) );
  INVX2 U14550 ( .A(n29191), .Y(n34338) );
  INVX1 U14551 ( .A(n31648), .Y(n25674) );
  INVX1 U14552 ( .A(n27020), .Y(n25675) );
  INVX1 U14553 ( .A(nc[9]), .Y(n25676) );
  INVX1 U14554 ( .A(n25676), .Y(n25677) );
  INVX1 U14555 ( .A(n25849), .Y(n25678) );
  INVX1 U14556 ( .A(n29423), .Y(n25679) );
  BUFX4 U14557 ( .A(n25641), .Y(n25680) );
  AND2X2 U14558 ( .A(n22988), .B(n25616), .Y(n25681) );
  INVX2 U14559 ( .A(n27913), .Y(n27915) );
  XNOR2X1 U14560 ( .A(n34390), .B(n21228), .Y(n34396) );
  INVX1 U14561 ( .A(n33123), .Y(n25682) );
  INVX1 U14562 ( .A(n25682), .Y(n25683) );
  INVX1 U14563 ( .A(n27903), .Y(n25684) );
  INVX4 U14564 ( .A(n25684), .Y(n25685) );
  INVX1 U14565 ( .A(net149876), .Y(net112194) );
  INVX1 U14566 ( .A(net111237), .Y(net112188) );
  AND2X2 U14567 ( .A(n32842), .B(n32841), .Y(n32843) );
  INVX1 U14568 ( .A(n29624), .Y(n25686) );
  INVX1 U14569 ( .A(net142728), .Y(net112181) );
  OAI21X1 U14570 ( .A(n27302), .B(n29465), .C(n27084), .Y(n25687) );
  XNOR2X1 U14571 ( .A(n33079), .B(n33099), .Y(n25699) );
  AND2X2 U14572 ( .A(oc[10]), .B(oc[8]), .Y(n29715) );
  OAI21X1 U14573 ( .A(n23139), .B(n25683), .C(n21363), .Y(n25690) );
  INVX1 U14574 ( .A(oc[0]), .Y(n25691) );
  INVX4 U14575 ( .A(n25691), .Y(n25692) );
  BUFX2 U14576 ( .A(n3159), .Y(n25693) );
  AND2X2 U14577 ( .A(n21142), .B(n23586), .Y(n25694) );
  INVX1 U14578 ( .A(n3200), .Y(n25695) );
  INVX1 U14579 ( .A(n25695), .Y(n25696) );
  MUX2X1 U14580 ( .B(n25699), .A(n25700), .S(n25730), .Y(n25698) );
  AND2X2 U14581 ( .A(n27178), .B(n25701), .Y(n25834) );
  AND2X2 U14582 ( .A(n34443), .B(n34360), .Y(n25701) );
  INVX2 U14583 ( .A(n25712), .Y(n25702) );
  INVX1 U14584 ( .A(n2246), .Y(n25703) );
  INVX1 U14585 ( .A(n25703), .Y(n25704) );
  INVX1 U14586 ( .A(n25688), .Y(n34442) );
  INVX1 U14587 ( .A(n32751), .Y(n25705) );
  INVX1 U14588 ( .A(n25715), .Y(n31917) );
  AND2X2 U14589 ( .A(n23086), .B(n33065), .Y(n25706) );
  INVX1 U14590 ( .A(n22966), .Y(n25707) );
  MUX2X1 U14591 ( .B(n28022), .A(n28021), .S(n29443), .Y(n28020) );
  MUX2X1 U14592 ( .B(n27991), .A(n27992), .S(n28221), .Y(n27990) );
  INVX4 U14593 ( .A(n29443), .Y(n28221) );
  INVX1 U14594 ( .A(oc[12]), .Y(n25708) );
  INVX4 U14595 ( .A(n25708), .Y(n25709) );
  INVX1 U14596 ( .A(n27903), .Y(n25710) );
  INVX4 U14597 ( .A(n25710), .Y(n25711) );
  INVX1 U14598 ( .A(oc[14]), .Y(n25712) );
  INVX1 U14599 ( .A(n25712), .Y(n25713) );
  NAND3X1 U14600 ( .A(net111332), .B(net115619), .C(net149940), .Y(n25716) );
  NAND3X1 U14601 ( .A(net95303), .B(n25727), .C(pLoc[0]), .Y(net111628) );
  INVX1 U14602 ( .A(nc[3]), .Y(n25717) );
  INVX1 U14603 ( .A(n25717), .Y(n25718) );
  INVX1 U14604 ( .A(n25689), .Y(n25719) );
  BUFX2 U14605 ( .A(n25687), .Y(n26164) );
  AND2X2 U14606 ( .A(n20977), .B(n27258), .Y(n25721) );
  MUX2X1 U14607 ( .B(n28129), .A(n28128), .S(n25732), .Y(n28127) );
  INVX1 U14608 ( .A(n25720), .Y(n25722) );
  INVX1 U14609 ( .A(n27253), .Y(n25723) );
  INVX1 U14610 ( .A(n25634), .Y(n25724) );
  AND2X2 U14611 ( .A(net110926), .B(net114252), .Y(n25727) );
  AND2X2 U14612 ( .A(n27903), .B(n22997), .Y(n25728) );
  MUX2X1 U14613 ( .B(grid[262]), .A(grid[256]), .S(net150787), .Y(n28180) );
  OAI21X1 U14614 ( .A(n22685), .B(n33097), .C(n33104), .Y(n25730) );
  MUX2X1 U14615 ( .B(grid[226]), .A(grid[220]), .S(net116755), .Y(n28182) );
  BUFX2 U14616 ( .A(n27319), .Y(n25731) );
  INVX4 U14617 ( .A(net106018), .Y(net53596) );
  INVX1 U14618 ( .A(n25744), .Y(n32514) );
  MUX2X1 U14619 ( .B(n34397), .A(n34396), .S(n34395), .Y(n25734) );
  INVX1 U14620 ( .A(n20992), .Y(n25735) );
  INVX1 U14621 ( .A(n29314), .Y(n25736) );
  INVX1 U14622 ( .A(n20993), .Y(n25737) );
  INVX1 U14623 ( .A(n20992), .Y(n25738) );
  INVX1 U14624 ( .A(n29314), .Y(n25739) );
  INVX1 U14625 ( .A(n20979), .Y(n25741) );
  INVX1 U14626 ( .A(n20988), .Y(n25742) );
  MUX2X1 U14627 ( .B(grid[247]), .A(grid[241]), .S(net150133), .Y(n27997) );
  AND2X2 U14628 ( .A(n23284), .B(n21106), .Y(n25743) );
  INVX2 U14629 ( .A(n25743), .Y(n32953) );
  NAND3X1 U14630 ( .A(n21360), .B(n25745), .C(n25746), .Y(n25744) );
  BUFX4 U14631 ( .A(n34426), .Y(n25748) );
  BUFX2 U14632 ( .A(n25483), .Y(n27178) );
  INVX1 U14633 ( .A(n22969), .Y(n25749) );
  INVX1 U14634 ( .A(n25194), .Y(n29993) );
  OAI21X1 U14635 ( .A(n34400), .B(n34405), .C(n34398), .Y(n25750) );
  BUFX2 U14636 ( .A(n3109), .Y(n25751) );
  MUX2X1 U14637 ( .B(n25405), .A(n25664), .S(n25681), .Y(n25752) );
  INVX4 U14638 ( .A(n26819), .Y(n33900) );
  MUX2X1 U14639 ( .B(grid[370]), .A(grid[364]), .S(net151633), .Y(n28161) );
  INVX1 U14640 ( .A(n20943), .Y(net110809) );
  INVX1 U14641 ( .A(n29557), .Y(n30050) );
  AND2X2 U14642 ( .A(n26070), .B(n25705), .Y(n25753) );
  INVX1 U14643 ( .A(alt14_net6192), .Y(net110686) );
  INVX1 U14644 ( .A(alt14_net6191), .Y(net110687) );
  INVX8 U14645 ( .A(n29383), .Y(n29381) );
  INVX1 U14646 ( .A(net110685), .Y(n4225) );
  INVX1 U14647 ( .A(net53623), .Y(net110421) );
  MUX2X1 U14648 ( .B(n28168), .A(n28167), .S(net105821), .Y(n28166) );
  NOR3X1 U14649 ( .A(n34230), .B(n21104), .C(n25825), .Y(n25754) );
  MUX2X1 U14650 ( .B(n28322), .A(n28321), .S(n26514), .Y(n28320) );
  AOI21X1 U14651 ( .A(n25329), .B(n33156), .C(n23426), .Y(n25755) );
  INVX2 U14652 ( .A(n25329), .Y(n33099) );
  INVX1 U14653 ( .A(n29247), .Y(n25757) );
  INVX1 U14654 ( .A(n29247), .Y(n25758) );
  INVX4 U14655 ( .A(n31885), .Y(n29247) );
  INVX1 U14656 ( .A(net151710), .Y(net89806) );
  INVX1 U14657 ( .A(n29511), .Y(n25760) );
  BUFX2 U14658 ( .A(n30652), .Y(n27172) );
  MUX2X1 U14659 ( .B(n25762), .A(n34248), .S(n23187), .Y(n25761) );
  INVX2 U14660 ( .A(n25761), .Y(n34249) );
  INVX1 U14661 ( .A(n23465), .Y(n25763) );
  AND2X2 U14662 ( .A(n22980), .B(n22994), .Y(n25764) );
  INVX1 U14663 ( .A(n21074), .Y(n29496) );
  INVX1 U14664 ( .A(n25671), .Y(n25765) );
  INVX1 U14665 ( .A(n34414), .Y(n25766) );
  OAI21X1 U14666 ( .A(n25688), .B(n26072), .C(n20969), .Y(n25768) );
  INVX1 U14667 ( .A(net94649), .Y(net110410) );
  INVX1 U14668 ( .A(net110410), .Y(net110411) );
  MUX2X1 U14669 ( .B(n21215), .A(grid[361]), .S(n33062), .Y(n27779) );
  INVX1 U14670 ( .A(n23092), .Y(n25769) );
  INVX1 U14671 ( .A(n25769), .Y(n25770) );
  BUFX2 U14672 ( .A(n29794), .Y(n25771) );
  INVX1 U14673 ( .A(n33429), .Y(n25773) );
  INVX4 U14674 ( .A(n25773), .Y(n25774) );
  INVX1 U14675 ( .A(n32742), .Y(n25775) );
  MUX2X1 U14676 ( .B(n27930), .A(n27945), .S(net109824), .Y(alt14_net6006) );
  INVX1 U14677 ( .A(net104479), .Y(net109824) );
  BUFX2 U14678 ( .A(n3154), .Y(n25776) );
  BUFX2 U14679 ( .A(n4226), .Y(net110320) );
  OR2X2 U14680 ( .A(n32616), .B(n32615), .Y(n32622) );
  MUX2X1 U14681 ( .B(grid[225]), .A(grid[219]), .S(net150133), .Y(n28122) );
  INVX1 U14682 ( .A(n21074), .Y(n25777) );
  INVX2 U14683 ( .A(n33085), .Y(n33154) );
  XNOR2X1 U14684 ( .A(n33074), .B(n33073), .Y(n33085) );
  AND2X2 U14685 ( .A(n27304), .B(n29697), .Y(n25779) );
  XNOR2X1 U14686 ( .A(n34393), .B(n25321), .Y(n25780) );
  INVX8 U14687 ( .A(n29461), .Y(n28607) );
  INVX1 U14688 ( .A(n29275), .Y(n25781) );
  INVX1 U14689 ( .A(n29275), .Y(n25782) );
  BUFX2 U14690 ( .A(n30665), .Y(n25783) );
  BUFX2 U14691 ( .A(n30665), .Y(n25784) );
  INVX1 U14692 ( .A(n25783), .Y(n25785) );
  INVX1 U14693 ( .A(n25783), .Y(n25786) );
  INVX1 U14694 ( .A(n25783), .Y(n25787) );
  INVX1 U14695 ( .A(n25783), .Y(n25788) );
  INVX1 U14696 ( .A(n25821), .Y(n25789) );
  INVX1 U14697 ( .A(n25821), .Y(n25790) );
  INVX1 U14698 ( .A(n25821), .Y(n25791) );
  INVX1 U14699 ( .A(n25821), .Y(n25792) );
  INVX1 U14700 ( .A(n25821), .Y(n25793) );
  INVX1 U14701 ( .A(n25821), .Y(n25794) );
  INVX1 U14702 ( .A(n25809), .Y(n25795) );
  INVX1 U14703 ( .A(n25821), .Y(n25796) );
  INVX1 U14704 ( .A(n25809), .Y(n25797) );
  INVX1 U14705 ( .A(n25784), .Y(n25798) );
  INVX1 U14706 ( .A(n25784), .Y(n25799) );
  INVX1 U14707 ( .A(n25784), .Y(n25800) );
  INVX1 U14708 ( .A(n25821), .Y(n25801) );
  INVX1 U14709 ( .A(n25783), .Y(n25802) );
  INVX1 U14710 ( .A(n25783), .Y(n25803) );
  INVX1 U14711 ( .A(n25783), .Y(n25804) );
  INVX1 U14712 ( .A(n25783), .Y(n25805) );
  INVX1 U14713 ( .A(n25781), .Y(n25806) );
  INVX1 U14714 ( .A(n25781), .Y(n25807) );
  INVX1 U14715 ( .A(n25781), .Y(n25808) );
  INVX1 U14716 ( .A(n25781), .Y(n25809) );
  INVX1 U14717 ( .A(n25806), .Y(n25810) );
  INVX1 U14718 ( .A(n25806), .Y(n25811) );
  INVX1 U14719 ( .A(n25806), .Y(n25812) );
  INVX1 U14720 ( .A(n25806), .Y(n25813) );
  INVX1 U14721 ( .A(n25806), .Y(n25814) );
  INVX1 U14722 ( .A(n25807), .Y(n25815) );
  INVX1 U14723 ( .A(n25807), .Y(n25816) );
  INVX1 U14724 ( .A(n25808), .Y(n25817) );
  INVX1 U14725 ( .A(n25808), .Y(n25818) );
  INVX1 U14726 ( .A(n25808), .Y(n25819) );
  INVX1 U14727 ( .A(n25809), .Y(n25820) );
  INVX1 U14728 ( .A(n25821), .Y(n25822) );
  INVX1 U14729 ( .A(n25821), .Y(n25823) );
  INVX1 U14730 ( .A(n25821), .Y(n25824) );
  INVX1 U14731 ( .A(n30665), .Y(n31907) );
  INVX1 U14732 ( .A(n34279), .Y(n25825) );
  INVX1 U14733 ( .A(n33154), .Y(n25826) );
  MUX2X1 U14734 ( .B(n34397), .A(n34396), .S(n34395), .Y(n25827) );
  OAI21X1 U14735 ( .A(n33120), .B(n25759), .C(n33119), .Y(n25828) );
  INVX8 U14736 ( .A(n28992), .Y(n27214) );
  AND2X2 U14737 ( .A(n9137), .B(n29381), .Y(n21794) );
  INVX4 U14738 ( .A(alt14_net96258), .Y(net105786) );
  INVX4 U14739 ( .A(net105786), .Y(net105788) );
  INVX1 U14740 ( .A(net151212), .Y(net95156) );
  INVX8 U14741 ( .A(n32773), .Y(n25830) );
  INVX1 U14742 ( .A(n27251), .Y(n25831) );
  INVX1 U14743 ( .A(n25756), .Y(n25832) );
  MUX2X1 U14744 ( .B(n28172), .A(n28187), .S(net109824), .Y(alt14_net6254) );
  AND2X2 U14745 ( .A(n29609), .B(n29608), .Y(n26069) );
  AND2X1 U14746 ( .A(n26896), .B(n29606), .Y(n29608) );
  MUX2X1 U14747 ( .B(n28160), .A(n28163), .S(alt14_net96304), .Y(n28174) );
  OAI21X1 U14748 ( .A(n25748), .B(n34425), .C(n34424), .Y(n25833) );
  INVX1 U14749 ( .A(n25834), .Y(n34302) );
  OR2X2 U14750 ( .A(n33006), .B(n33005), .Y(n33013) );
  INVX2 U14751 ( .A(n27251), .Y(n25839) );
  INVX1 U14752 ( .A(n22673), .Y(n25836) );
  INVX1 U14753 ( .A(n34352), .Y(n25837) );
  INVX1 U14754 ( .A(n25837), .Y(n25838) );
  INVX1 U14755 ( .A(n29513), .Y(n25840) );
  OR2X2 U14756 ( .A(n21057), .B(n29353), .Y(n30642) );
  INVX8 U14757 ( .A(n29353), .Y(n29352) );
  INVX1 U14758 ( .A(n29633), .Y(n25841) );
  BUFX4 U14759 ( .A(n2249), .Y(n28993) );
  INVX1 U14760 ( .A(n31493), .Y(n25842) );
  AND2X2 U14761 ( .A(n25466), .B(n31482), .Y(n25843) );
  INVX1 U14762 ( .A(n25852), .Y(n25844) );
  AND2X2 U14763 ( .A(n23644), .B(n25196), .Y(n25845) );
  INVX1 U14764 ( .A(n25845), .Y(n33112) );
  INVX1 U14765 ( .A(n21196), .Y(n25846) );
  NAND3X1 U14766 ( .A(n29503), .B(n21058), .C(n23140), .Y(n25847) );
  INVX2 U14767 ( .A(alt5_net95668), .Y(alt5_net95666) );
  INVX2 U14768 ( .A(alt5_net95668), .Y(alt5_net95664) );
  AND2X2 U14769 ( .A(states[0]), .B(n29603), .Y(net109585) );
  INVX1 U14770 ( .A(alt14_net6005), .Y(net108805) );
  INVX1 U14771 ( .A(n34383), .Y(n25851) );
  INVX2 U14772 ( .A(n34382), .Y(n34383) );
  INVX1 U14773 ( .A(net143109), .Y(net109485) );
  BUFX2 U14774 ( .A(n4224), .Y(net109469) );
  INVX1 U14775 ( .A(n25678), .Y(n25852) );
  INVX2 U14776 ( .A(n29248), .Y(n25853) );
  INVX8 U14777 ( .A(n25853), .Y(n25854) );
  INVX1 U14778 ( .A(n31885), .Y(n29248) );
  INVX1 U14779 ( .A(net138174), .Y(net109440) );
  MUX2X1 U14780 ( .B(n25204), .A(n24324), .S(n33071), .Y(n33074) );
  INVX1 U14781 ( .A(n29247), .Y(n25856) );
  INVX1 U14782 ( .A(n29247), .Y(n25857) );
  INVX1 U14783 ( .A(n34414), .Y(n25858) );
  XNOR2X1 U14784 ( .A(n23104), .B(n34317), .Y(n34315) );
  XNOR2X1 U14785 ( .A(n25827), .B(n34400), .Y(n25860) );
  INVX1 U14786 ( .A(n25734), .Y(n34404) );
  INVX1 U14787 ( .A(n34420), .Y(n25861) );
  AND2X2 U14788 ( .A(n34374), .B(n34372), .Y(n25863) );
  INVX1 U14789 ( .A(n25863), .Y(n34391) );
  INVX1 U14790 ( .A(alt14_net6006), .Y(net108804) );
  XNOR2X1 U14791 ( .A(n27913), .B(n34385), .Y(n25864) );
  INVX2 U14792 ( .A(n25864), .Y(n34378) );
  INVX8 U14793 ( .A(n25839), .Y(n27913) );
  INVX1 U14794 ( .A(n23201), .Y(n25865) );
  INVX1 U14795 ( .A(n29273), .Y(n25866) );
  BUFX2 U14796 ( .A(n29273), .Y(n25867) );
  BUFX2 U14797 ( .A(n29273), .Y(n25868) );
  BUFX2 U14798 ( .A(n29273), .Y(n25869) );
  INVX1 U14799 ( .A(n25867), .Y(n25870) );
  INVX1 U14800 ( .A(n25868), .Y(n25871) );
  INVX1 U14801 ( .A(n25869), .Y(n25872) );
  BUFX2 U14802 ( .A(n25413), .Y(n25873) );
  BUFX2 U14803 ( .A(n25413), .Y(n25874) );
  BUFX2 U14804 ( .A(n25413), .Y(n25875) );
  INVX1 U14805 ( .A(n25873), .Y(n25876) );
  INVX1 U14806 ( .A(n25873), .Y(n25877) );
  INVX1 U14807 ( .A(n25873), .Y(n25878) );
  INVX1 U14808 ( .A(n25873), .Y(n25879) );
  INVX1 U14809 ( .A(n25874), .Y(n25880) );
  INVX1 U14810 ( .A(n25874), .Y(n25881) );
  INVX1 U14811 ( .A(n25874), .Y(n25882) );
  INVX1 U14812 ( .A(n25874), .Y(n25883) );
  INVX1 U14813 ( .A(n25875), .Y(n25884) );
  INVX1 U14814 ( .A(n25875), .Y(n25885) );
  INVX1 U14815 ( .A(n25875), .Y(n25886) );
  INVX1 U14816 ( .A(n25875), .Y(n25887) );
  BUFX2 U14817 ( .A(n29272), .Y(n25888) );
  BUFX2 U14818 ( .A(n29272), .Y(n25889) );
  BUFX2 U14819 ( .A(n29272), .Y(n25890) );
  INVX1 U14820 ( .A(n25888), .Y(n25891) );
  INVX1 U14821 ( .A(n25888), .Y(n25892) );
  INVX1 U14822 ( .A(n25888), .Y(n25893) );
  INVX1 U14823 ( .A(n25888), .Y(n25894) );
  INVX1 U14824 ( .A(n25889), .Y(n25895) );
  INVX1 U14825 ( .A(n25889), .Y(n25896) );
  INVX1 U14826 ( .A(n25889), .Y(n25897) );
  INVX1 U14827 ( .A(n25889), .Y(n25898) );
  INVX1 U14828 ( .A(n25890), .Y(n25899) );
  INVX1 U14829 ( .A(n25890), .Y(n25900) );
  INVX1 U14830 ( .A(n25890), .Y(n25901) );
  INVX1 U14831 ( .A(n25890), .Y(n25902) );
  INVX1 U14832 ( .A(n25414), .Y(n25903) );
  INVX1 U14833 ( .A(n25414), .Y(n25904) );
  INVX1 U14834 ( .A(n25414), .Y(n25905) );
  INVX1 U14835 ( .A(n25414), .Y(n25906) );
  INVX1 U14836 ( .A(n25903), .Y(n25907) );
  INVX1 U14837 ( .A(n25903), .Y(n25908) );
  INVX1 U14838 ( .A(n25903), .Y(n25909) );
  INVX1 U14839 ( .A(n25903), .Y(n25910) );
  INVX1 U14840 ( .A(n25904), .Y(n25911) );
  INVX1 U14841 ( .A(n25904), .Y(n25912) );
  INVX1 U14842 ( .A(n25904), .Y(n25913) );
  INVX1 U14843 ( .A(n25904), .Y(n25914) );
  INVX1 U14844 ( .A(n25905), .Y(n25915) );
  INVX1 U14845 ( .A(n25905), .Y(n25916) );
  INVX1 U14846 ( .A(n25905), .Y(n25917) );
  INVX1 U14847 ( .A(n25905), .Y(n25918) );
  INVX1 U14848 ( .A(n25906), .Y(n25919) );
  INVX1 U14849 ( .A(n25906), .Y(n25920) );
  INVX1 U14850 ( .A(n25906), .Y(n25921) );
  INVX1 U14851 ( .A(n25906), .Y(n25922) );
  INVX1 U14852 ( .A(n25866), .Y(n25923) );
  INVX1 U14853 ( .A(n25866), .Y(n25924) );
  INVX1 U14854 ( .A(n25923), .Y(n25925) );
  INVX1 U14855 ( .A(n25923), .Y(n25926) );
  INVX1 U14856 ( .A(n25923), .Y(n25927) );
  INVX1 U14857 ( .A(n25923), .Y(n25928) );
  INVX1 U14858 ( .A(n25924), .Y(n25929) );
  INVX1 U14859 ( .A(n25924), .Y(n25930) );
  INVX1 U14860 ( .A(n25924), .Y(n25931) );
  INVX1 U14861 ( .A(net94647), .Y(net109176) );
  INVX1 U14862 ( .A(n29276), .Y(n25932) );
  INVX1 U14863 ( .A(n29276), .Y(n25933) );
  BUFX2 U14864 ( .A(n30686), .Y(n25934) );
  BUFX2 U14865 ( .A(n30686), .Y(n25935) );
  BUFX2 U14866 ( .A(n30686), .Y(n25936) );
  INVX1 U14867 ( .A(n25934), .Y(n25937) );
  INVX1 U14868 ( .A(n25934), .Y(n25938) );
  INVX1 U14869 ( .A(n25934), .Y(n25939) );
  INVX1 U14870 ( .A(n25934), .Y(n25940) );
  INVX1 U14871 ( .A(n21092), .Y(n25941) );
  INVX1 U14872 ( .A(n25935), .Y(n25942) );
  INVX1 U14873 ( .A(n25935), .Y(n25943) );
  INVX1 U14874 ( .A(n25935), .Y(n25944) );
  INVX1 U14875 ( .A(n25935), .Y(n25945) );
  INVX1 U14876 ( .A(n25935), .Y(n25946) );
  INVX1 U14877 ( .A(n21092), .Y(n25947) );
  INVX1 U14878 ( .A(n21092), .Y(n25948) );
  INVX1 U14879 ( .A(n25936), .Y(n25949) );
  INVX1 U14880 ( .A(n25936), .Y(n25950) );
  INVX1 U14881 ( .A(n25936), .Y(n25951) );
  INVX1 U14882 ( .A(n25936), .Y(n25952) );
  INVX1 U14883 ( .A(n25936), .Y(n25953) );
  INVX1 U14884 ( .A(n25934), .Y(n25954) );
  INVX1 U14885 ( .A(n25934), .Y(n25955) );
  INVX1 U14886 ( .A(n25932), .Y(n25956) );
  INVX1 U14887 ( .A(n25932), .Y(n25957) );
  INVX1 U14888 ( .A(n25932), .Y(n25958) );
  INVX1 U14889 ( .A(n25956), .Y(n25959) );
  INVX1 U14890 ( .A(n25956), .Y(n25960) );
  INVX1 U14891 ( .A(n25956), .Y(n25961) );
  INVX1 U14892 ( .A(n25957), .Y(n25962) );
  INVX1 U14893 ( .A(n25957), .Y(n25963) );
  INVX1 U14894 ( .A(n25957), .Y(n25964) );
  INVX1 U14895 ( .A(n25958), .Y(n25965) );
  INVX1 U14896 ( .A(n25958), .Y(n25966) );
  INVX1 U14897 ( .A(n25958), .Y(n25967) );
  INVX1 U14898 ( .A(n25972), .Y(n25968) );
  INVX1 U14899 ( .A(n25971), .Y(n25969) );
  INVX1 U14900 ( .A(n21092), .Y(n25970) );
  INVX1 U14901 ( .A(n25933), .Y(n25971) );
  INVX1 U14902 ( .A(n25933), .Y(n25972) );
  INVX1 U14903 ( .A(n25933), .Y(n25973) );
  INVX1 U14904 ( .A(n25971), .Y(n25974) );
  INVX1 U14905 ( .A(n25972), .Y(n25975) );
  INVX1 U14906 ( .A(n25972), .Y(n25976) );
  INVX1 U14907 ( .A(n25973), .Y(n25977) );
  INVX1 U14908 ( .A(n25973), .Y(n25978) );
  INVX1 U14909 ( .A(n25973), .Y(n25979) );
  INVX1 U14910 ( .A(n30686), .Y(n31908) );
  INVX1 U14911 ( .A(n29250), .Y(n25980) );
  BUFX2 U14912 ( .A(n29249), .Y(n25981) );
  BUFX2 U14913 ( .A(n29249), .Y(n25982) );
  BUFX2 U14914 ( .A(n29250), .Y(n25983) );
  INVX1 U14915 ( .A(n25981), .Y(n25984) );
  INVX1 U14916 ( .A(n25981), .Y(n25985) );
  INVX1 U14917 ( .A(n25981), .Y(n25986) );
  INVX1 U14918 ( .A(n25981), .Y(n25987) );
  INVX1 U14919 ( .A(n25982), .Y(n25988) );
  INVX1 U14920 ( .A(n25982), .Y(n25989) );
  INVX1 U14921 ( .A(n25982), .Y(n25990) );
  INVX1 U14922 ( .A(n25982), .Y(n25991) );
  INVX1 U14923 ( .A(n25983), .Y(n25992) );
  INVX1 U14924 ( .A(n25983), .Y(n25993) );
  INVX1 U14925 ( .A(n25983), .Y(n25994) );
  INVX1 U14926 ( .A(n25983), .Y(n25995) );
  BUFX2 U14927 ( .A(n29252), .Y(n25996) );
  INVX1 U14928 ( .A(n25996), .Y(n25997) );
  INVX1 U14929 ( .A(n25996), .Y(n25998) );
  INVX1 U14930 ( .A(n25996), .Y(n25999) );
  INVX1 U14931 ( .A(n25996), .Y(n26000) );
  BUFX2 U14932 ( .A(n21000), .Y(n26001) );
  BUFX2 U14933 ( .A(n21000), .Y(n26002) );
  BUFX2 U14934 ( .A(n21000), .Y(n26003) );
  INVX1 U14935 ( .A(n26001), .Y(n26004) );
  INVX1 U14936 ( .A(n26001), .Y(n26005) );
  INVX1 U14937 ( .A(n26001), .Y(n26006) );
  INVX1 U14938 ( .A(n26001), .Y(n26007) );
  INVX1 U14939 ( .A(n26002), .Y(n26008) );
  INVX1 U14940 ( .A(n26002), .Y(n26009) );
  INVX1 U14941 ( .A(n26002), .Y(n26010) );
  INVX1 U14942 ( .A(n26002), .Y(n26011) );
  INVX1 U14943 ( .A(n26003), .Y(n26012) );
  INVX1 U14944 ( .A(n26003), .Y(n26013) );
  INVX1 U14945 ( .A(n26003), .Y(n26014) );
  INVX1 U14946 ( .A(n26003), .Y(n26015) );
  INVX1 U14947 ( .A(n25412), .Y(n26016) );
  INVX1 U14948 ( .A(n25412), .Y(n26017) );
  INVX1 U14949 ( .A(n25412), .Y(n26018) );
  INVX1 U14950 ( .A(n25412), .Y(n26019) );
  INVX1 U14951 ( .A(n26016), .Y(n26020) );
  INVX1 U14952 ( .A(n26016), .Y(n26021) );
  INVX1 U14953 ( .A(n26017), .Y(n26022) );
  INVX1 U14954 ( .A(n26017), .Y(n26023) );
  INVX1 U14955 ( .A(n26017), .Y(n26024) );
  INVX1 U14956 ( .A(n26017), .Y(n26025) );
  INVX1 U14957 ( .A(n26018), .Y(n26026) );
  INVX1 U14958 ( .A(n26018), .Y(n26027) );
  INVX1 U14959 ( .A(n26018), .Y(n26028) );
  INVX1 U14960 ( .A(n26018), .Y(n26029) );
  INVX1 U14961 ( .A(n26019), .Y(n26030) );
  INVX1 U14962 ( .A(n26019), .Y(n26031) );
  INVX1 U14963 ( .A(n26019), .Y(n26032) );
  INVX1 U14964 ( .A(n26019), .Y(n26033) );
  INVX1 U14965 ( .A(n25980), .Y(n26034) );
  INVX1 U14966 ( .A(n25980), .Y(n26035) );
  INVX1 U14967 ( .A(n26034), .Y(n26036) );
  INVX1 U14968 ( .A(n26034), .Y(n26037) );
  INVX1 U14969 ( .A(n26034), .Y(n26038) );
  INVX1 U14970 ( .A(n26034), .Y(n26039) );
  INVX1 U14971 ( .A(n26035), .Y(n26040) );
  INVX1 U14972 ( .A(n26035), .Y(n26041) );
  INVX1 U14973 ( .A(n26035), .Y(n26042) );
  XNOR2X1 U14974 ( .A(n34304), .B(n26044), .Y(n26043) );
  AND2X2 U14975 ( .A(n21988), .B(n25629), .Y(n26044) );
  INVX1 U14976 ( .A(n29383), .Y(n29379) );
  INVX1 U14977 ( .A(n33144), .Y(n26045) );
  AND2X2 U14978 ( .A(n34292), .B(n34356), .Y(n26046) );
  MUX2X1 U14979 ( .B(n27792), .A(n27791), .S(n25611), .Y(n27790) );
  OR2X2 U14980 ( .A(n25768), .B(T[5]), .Y(n33104) );
  INVX1 U14981 ( .A(n22964), .Y(n26047) );
  INVX1 U14982 ( .A(n26047), .Y(n26048) );
  AND2X2 U14983 ( .A(n23001), .B(n34298), .Y(n26049) );
  NOR3X1 U14984 ( .A(n26051), .B(alt5_net95668), .C(n29178), .Y(n26050) );
  BUFX2 U14985 ( .A(oc[26]), .Y(n26052) );
  INVX1 U14986 ( .A(n26045), .Y(n26053) );
  INVX1 U14987 ( .A(n34362), .Y(n26054) );
  INVX1 U14988 ( .A(n25779), .Y(n26056) );
  INVX1 U14989 ( .A(net109585), .Y(net108653) );
  OAI21X1 U14990 ( .A(n25838), .B(n34351), .C(n27158), .Y(n26058) );
  INVX1 U14991 ( .A(net94645), .Y(net108619) );
  INVX1 U14992 ( .A(n34424), .Y(n26059) );
  BUFX2 U14993 ( .A(n23467), .Y(n26060) );
  BUFX2 U14994 ( .A(n22673), .Y(n26062) );
  INVX1 U14995 ( .A(n22964), .Y(n29466) );
  INVX1 U14996 ( .A(net111332), .Y(n4125) );
  INVX1 U14997 ( .A(n20808), .Y(n26064) );
  INVX1 U14998 ( .A(n26064), .Y(n26065) );
  INVX1 U14999 ( .A(oc[19]), .Y(n26067) );
  INVX4 U15000 ( .A(n26067), .Y(n26068) );
  INVX2 U15001 ( .A(oc[31]), .Y(n29725) );
  INVX1 U15002 ( .A(n32472), .Y(n26071) );
  AND2X2 U15003 ( .A(n9134), .B(n29381), .Y(n21791) );
  AND2X2 U15004 ( .A(n33049), .B(n33050), .Y(n29193) );
  INVX8 U15005 ( .A(n27913), .Y(n27914) );
  AND2X2 U15006 ( .A(n32511), .B(n32510), .Y(n32512) );
  INVX4 U15007 ( .A(n34315), .Y(n34434) );
  AND2X2 U15008 ( .A(n20977), .B(n29679), .Y(n27264) );
  AND2X2 U15009 ( .A(n27310), .B(n21186), .Y(n27266) );
  INVX1 U15010 ( .A(n2252), .Y(n26073) );
  INVX1 U15011 ( .A(n29183), .Y(n26074) );
  INVX1 U15012 ( .A(n29180), .Y(n26075) );
  INVX1 U15013 ( .A(n29181), .Y(n26076) );
  INVX8 U15014 ( .A(n29179), .Y(n29182) );
  INVX2 U15015 ( .A(n29179), .Y(n29181) );
  INVX4 U15016 ( .A(n2252), .Y(n29179) );
  AND2X2 U15017 ( .A(n27258), .B(n21183), .Y(n27306) );
  AND2X2 U15018 ( .A(n27310), .B(n21183), .Y(n27305) );
  AND2X2 U15019 ( .A(n29509), .B(n29477), .Y(n27256) );
  AND2X2 U15020 ( .A(n23290), .B(n29331), .Y(n27216) );
  AND2X2 U15021 ( .A(n23285), .B(n25724), .Y(n27217) );
  AND2X2 U15022 ( .A(n22992), .B(n25849), .Y(n27295) );
  INVX4 U15023 ( .A(n27190), .Y(n33806) );
  AND2X2 U15024 ( .A(n27244), .B(net150133), .Y(n27222) );
  INVX1 U15025 ( .A(n26484), .Y(n26079) );
  INVX1 U15026 ( .A(n26446), .Y(n26080) );
  INVX1 U15027 ( .A(n21097), .Y(n26081) );
  INVX1 U15028 ( .A(n26517), .Y(n26082) );
  INVX1 U15029 ( .A(n26484), .Y(n26083) );
  INVX1 U15030 ( .A(n21163), .Y(n26085) );
  INVX1 U15031 ( .A(n26445), .Y(n26086) );
  INVX1 U15032 ( .A(n26445), .Y(n26088) );
  INVX1 U15033 ( .A(n26445), .Y(n26089) );
  INVX1 U15034 ( .A(n26445), .Y(n26091) );
  INVX1 U15035 ( .A(n26445), .Y(n26092) );
  INVX1 U15036 ( .A(n26445), .Y(n26093) );
  INVX1 U15037 ( .A(n28595), .Y(n26094) );
  INVX1 U15038 ( .A(n28595), .Y(n26095) );
  INVX1 U15039 ( .A(n26445), .Y(n26097) );
  INVX1 U15040 ( .A(n28595), .Y(n26098) );
  INVX1 U15041 ( .A(n28595), .Y(n26099) );
  INVX1 U15042 ( .A(n28595), .Y(n26100) );
  INVX1 U15043 ( .A(n26484), .Y(n26101) );
  INVX1 U15044 ( .A(n28595), .Y(n26103) );
  INVX1 U15045 ( .A(n26517), .Y(n26104) );
  INVX1 U15046 ( .A(n21163), .Y(n26105) );
  INVX1 U15047 ( .A(n26517), .Y(n26106) );
  INVX1 U15048 ( .A(n28595), .Y(n26107) );
  INVX1 U15049 ( .A(n26517), .Y(n26108) );
  INVX1 U15050 ( .A(n28595), .Y(n26109) );
  INVX1 U15051 ( .A(n28595), .Y(n26110) );
  INVX1 U15052 ( .A(n28595), .Y(n26111) );
  INVX1 U15053 ( .A(n28595), .Y(n26112) );
  INVX1 U15054 ( .A(n26445), .Y(n26113) );
  INVX1 U15055 ( .A(n26484), .Y(n26114) );
  INVX1 U15056 ( .A(n28595), .Y(n26117) );
  INVX1 U15057 ( .A(n26517), .Y(n26118) );
  INVX1 U15058 ( .A(n26445), .Y(n26119) );
  INVX1 U15059 ( .A(n26445), .Y(n26120) );
  INVX1 U15060 ( .A(n21163), .Y(n26123) );
  INVX1 U15061 ( .A(n21163), .Y(n26124) );
  INVX1 U15062 ( .A(n26517), .Y(n26125) );
  INVX1 U15063 ( .A(n26484), .Y(n26126) );
  INVX1 U15064 ( .A(n21163), .Y(n26128) );
  INVX1 U15065 ( .A(n21163), .Y(n26129) );
  INVX1 U15066 ( .A(n28594), .Y(n26130) );
  INVX1 U15067 ( .A(n26516), .Y(n26131) );
  INVX1 U15068 ( .A(n21163), .Y(n26132) );
  INVX1 U15069 ( .A(n26517), .Y(n26133) );
  INVX1 U15070 ( .A(n26446), .Y(n26134) );
  INVX1 U15071 ( .A(n26446), .Y(n26135) );
  INVX1 U15072 ( .A(n26446), .Y(n26136) );
  INVX1 U15073 ( .A(n26484), .Y(n26137) );
  INVX1 U15074 ( .A(n21163), .Y(n26138) );
  INVX1 U15075 ( .A(n26484), .Y(n26140) );
  INVX1 U15076 ( .A(n26445), .Y(n26141) );
  INVX1 U15077 ( .A(n21163), .Y(n26142) );
  INVX1 U15078 ( .A(n26517), .Y(n26143) );
  INVX1 U15079 ( .A(n26517), .Y(n26144) );
  INVX1 U15080 ( .A(n26517), .Y(n26145) );
  INVX1 U15081 ( .A(n21163), .Y(n26147) );
  INVX1 U15082 ( .A(n21163), .Y(n26149) );
  INVX1 U15083 ( .A(n21163), .Y(n26150) );
  INVX1 U15084 ( .A(n21163), .Y(n26151) );
  INVX1 U15085 ( .A(n26516), .Y(n26152) );
  INVX1 U15086 ( .A(n26517), .Y(n26153) );
  INVX1 U15087 ( .A(n21097), .Y(n26154) );
  INVX1 U15088 ( .A(n21090), .Y(n26155) );
  INVX1 U15089 ( .A(n21090), .Y(n26156) );
  INVX1 U15090 ( .A(n26516), .Y(n26157) );
  INVX1 U15091 ( .A(n26516), .Y(n26158) );
  INVX1 U15092 ( .A(n21091), .Y(n26159) );
  INVX1 U15093 ( .A(n21091), .Y(n26160) );
  INVX1 U15094 ( .A(n21090), .Y(n26161) );
  INVX4 U15095 ( .A(n28598), .Y(n26517) );
  INVX1 U15096 ( .A(n26259), .Y(n26165) );
  INVX1 U15097 ( .A(n26259), .Y(n26166) );
  INVX1 U15098 ( .A(n26259), .Y(n26167) );
  INVX1 U15099 ( .A(n26260), .Y(n26168) );
  INVX1 U15100 ( .A(n26260), .Y(n26169) );
  INVX1 U15101 ( .A(n26259), .Y(n26170) );
  INVX1 U15102 ( .A(n26260), .Y(n26171) );
  BUFX4 U15103 ( .A(n26165), .Y(n26172) );
  BUFX4 U15104 ( .A(n26166), .Y(n26173) );
  BUFX4 U15105 ( .A(n26167), .Y(n26174) );
  INVX1 U15106 ( .A(n28987), .Y(n26179) );
  INVX1 U15107 ( .A(n28987), .Y(n26180) );
  INVX1 U15108 ( .A(n28987), .Y(n26181) );
  BUFX2 U15109 ( .A(n26179), .Y(n26182) );
  BUFX2 U15110 ( .A(n26180), .Y(n26183) );
  BUFX2 U15111 ( .A(n26181), .Y(n26184) );
  BUFX2 U15112 ( .A(n26180), .Y(n26185) );
  BUFX2 U15113 ( .A(n26180), .Y(n26186) );
  BUFX2 U15114 ( .A(n26181), .Y(n26187) );
  BUFX2 U15115 ( .A(n26181), .Y(n26188) );
  INVX1 U15116 ( .A(n28984), .Y(n26189) );
  INVX1 U15117 ( .A(n28984), .Y(n26190) );
  INVX1 U15118 ( .A(n28984), .Y(n26191) );
  INVX1 U15119 ( .A(n28984), .Y(n26192) );
  INVX1 U15120 ( .A(n28984), .Y(n26193) );
  INVX1 U15121 ( .A(n28984), .Y(n26194) );
  INVX1 U15122 ( .A(n28984), .Y(n26195) );
  BUFX4 U15123 ( .A(n26189), .Y(n26196) );
  BUFX4 U15124 ( .A(n26190), .Y(n26197) );
  BUFX4 U15125 ( .A(n26191), .Y(n26198) );
  BUFX4 U15126 ( .A(n26192), .Y(n26199) );
  BUFX4 U15127 ( .A(n26193), .Y(n26200) );
  BUFX4 U15128 ( .A(n26194), .Y(n26201) );
  BUFX4 U15129 ( .A(n26195), .Y(n26202) );
  INVX1 U15130 ( .A(n28983), .Y(n26203) );
  INVX1 U15131 ( .A(n28983), .Y(n26204) );
  INVX1 U15132 ( .A(n28983), .Y(n26205) );
  INVX1 U15133 ( .A(n28983), .Y(n26206) );
  INVX1 U15134 ( .A(n28983), .Y(n26207) );
  INVX1 U15135 ( .A(n28983), .Y(n26208) );
  INVX1 U15136 ( .A(n28983), .Y(n26209) );
  BUFX4 U15137 ( .A(n26203), .Y(n26210) );
  BUFX2 U15138 ( .A(n26204), .Y(n26211) );
  BUFX2 U15139 ( .A(n26205), .Y(n26212) );
  BUFX4 U15140 ( .A(n26206), .Y(n26213) );
  BUFX4 U15141 ( .A(n26207), .Y(n26214) );
  BUFX4 U15142 ( .A(n26208), .Y(n26215) );
  BUFX4 U15143 ( .A(n26209), .Y(n26216) );
  INVX1 U15144 ( .A(n28982), .Y(n26217) );
  INVX1 U15145 ( .A(n28982), .Y(n26218) );
  INVX1 U15146 ( .A(n28982), .Y(n26219) );
  INVX1 U15147 ( .A(n28982), .Y(n26220) );
  INVX1 U15148 ( .A(n28982), .Y(n26221) );
  INVX1 U15149 ( .A(n28982), .Y(n26222) );
  INVX1 U15150 ( .A(n28982), .Y(n26223) );
  BUFX4 U15151 ( .A(n26217), .Y(n26224) );
  BUFX4 U15152 ( .A(n26218), .Y(n26225) );
  BUFX4 U15153 ( .A(n26219), .Y(n26226) );
  BUFX4 U15154 ( .A(n26220), .Y(n26227) );
  BUFX4 U15155 ( .A(n26221), .Y(n26228) );
  BUFX4 U15156 ( .A(n26222), .Y(n26229) );
  BUFX4 U15157 ( .A(n26223), .Y(n26230) );
  INVX1 U15158 ( .A(n28985), .Y(n26231) );
  INVX1 U15159 ( .A(n28985), .Y(n26232) );
  INVX1 U15160 ( .A(n28985), .Y(n26233) );
  INVX1 U15161 ( .A(n28985), .Y(n26234) );
  INVX1 U15162 ( .A(n28985), .Y(n26235) );
  INVX1 U15163 ( .A(n28985), .Y(n26236) );
  INVX1 U15164 ( .A(n28985), .Y(n26237) );
  BUFX4 U15165 ( .A(n26231), .Y(n26238) );
  BUFX4 U15166 ( .A(n26232), .Y(n26239) );
  BUFX4 U15167 ( .A(n26233), .Y(n26240) );
  BUFX4 U15168 ( .A(n26234), .Y(n26241) );
  BUFX4 U15169 ( .A(n26235), .Y(n26242) );
  BUFX4 U15170 ( .A(n26236), .Y(n26243) );
  BUFX4 U15171 ( .A(n26237), .Y(n26244) );
  INVX1 U15172 ( .A(n28986), .Y(n26245) );
  INVX1 U15173 ( .A(n28986), .Y(n26246) );
  INVX1 U15174 ( .A(n28986), .Y(n26247) );
  INVX1 U15175 ( .A(n28986), .Y(n26248) );
  INVX1 U15176 ( .A(n28986), .Y(n26249) );
  INVX1 U15177 ( .A(n28986), .Y(n26250) );
  INVX1 U15178 ( .A(n28986), .Y(n26251) );
  BUFX4 U15179 ( .A(n26245), .Y(n26252) );
  BUFX4 U15180 ( .A(n26246), .Y(n26253) );
  BUFX4 U15181 ( .A(n26247), .Y(n26254) );
  BUFX4 U15182 ( .A(n26248), .Y(n26255) );
  BUFX4 U15183 ( .A(n26249), .Y(n26256) );
  BUFX4 U15184 ( .A(n26250), .Y(n26257) );
  BUFX4 U15185 ( .A(n26251), .Y(n26258) );
  INVX2 U15186 ( .A(n2245), .Y(n26259) );
  INVX2 U15187 ( .A(n2245), .Y(n26260) );
  INVX4 U15188 ( .A(n26259), .Y(n26261) );
  INVX4 U15189 ( .A(n26259), .Y(n26262) );
  INVX4 U15190 ( .A(n26260), .Y(n26263) );
  INVX4 U15191 ( .A(n26260), .Y(n26264) );
  INVX4 U15192 ( .A(n26260), .Y(n26265) );
  INVX2 U15193 ( .A(n26259), .Y(n26266) );
  INVX2 U15194 ( .A(n26259), .Y(n26267) );
  OR2X2 U15195 ( .A(n8034), .B(n8035), .Y(n30638) );
  AND2X2 U15196 ( .A(n30186), .B(n30281), .Y(n27258) );
  INVX1 U15197 ( .A(n22968), .Y(n34498) );
  INVX4 U15198 ( .A(n27102), .Y(n33875) );
  AND2X2 U15199 ( .A(n23282), .B(n29330), .Y(n27232) );
  AND2X2 U15200 ( .A(n32700), .B(n32699), .Y(n32701) );
  INVX1 U15201 ( .A(n21207), .Y(n26270) );
  INVX1 U15202 ( .A(n26270), .Y(n26271) );
  INVX1 U15203 ( .A(n32042), .Y(n26273) );
  INVX1 U15204 ( .A(n26273), .Y(n26274) );
  INVX1 U15205 ( .A(n25205), .Y(n26275) );
  INVX1 U15206 ( .A(n22971), .Y(n26276) );
  INVX1 U15207 ( .A(n26276), .Y(n26277) );
  INVX1 U15208 ( .A(n26278), .Y(n26279) );
  INVX1 U15209 ( .A(n26278), .Y(n26280) );
  INVX1 U15210 ( .A(n29230), .Y(n26281) );
  INVX1 U15211 ( .A(n26300), .Y(n26282) );
  INVX1 U15212 ( .A(n26300), .Y(n26283) );
  INVX1 U15213 ( .A(n26289), .Y(n26284) );
  INVX1 U15214 ( .A(n26289), .Y(n26285) );
  INVX1 U15215 ( .A(n26280), .Y(n26286) );
  INVX1 U15216 ( .A(n26295), .Y(n26287) );
  INVX1 U15217 ( .A(n29229), .Y(n26288) );
  INVX1 U15218 ( .A(n29229), .Y(n26289) );
  INVX1 U15219 ( .A(n26289), .Y(n26290) );
  INVX1 U15220 ( .A(n26288), .Y(n26291) );
  INVX1 U15221 ( .A(n22971), .Y(n26292) );
  INVX1 U15222 ( .A(n26276), .Y(n26295) );
  INVX1 U15223 ( .A(n26294), .Y(n26296) );
  INVX1 U15224 ( .A(n26294), .Y(n26297) );
  INVX1 U15225 ( .A(n26277), .Y(n26298) );
  INVX1 U15226 ( .A(n26301), .Y(n26299) );
  INVX1 U15227 ( .A(n29230), .Y(n26300) );
  INVX1 U15228 ( .A(n26292), .Y(n26301) );
  INVX1 U15229 ( .A(n26300), .Y(n26302) );
  INVX1 U15230 ( .A(n26301), .Y(n26303) );
  INVX1 U15231 ( .A(n29195), .Y(n29229) );
  AND2X2 U15232 ( .A(n32797), .B(n32796), .Y(n32798) );
  INVX1 U15233 ( .A(net117301), .Y(net107063) );
  INVX1 U15234 ( .A(net142728), .Y(net107074) );
  INVX1 U15235 ( .A(net142728), .Y(net107076) );
  INVX1 U15236 ( .A(net107074), .Y(net107078) );
  INVX1 U15237 ( .A(net151812), .Y(net107082) );
  INVX1 U15238 ( .A(net147983), .Y(net107088) );
  INVX1 U15239 ( .A(net112181), .Y(net107090) );
  INVX1 U15240 ( .A(net107076), .Y(net107091) );
  BUFX4 U15241 ( .A(n8052), .Y(n26304) );
  INVX1 U15242 ( .A(n29253), .Y(n26305) );
  INVX1 U15243 ( .A(n29253), .Y(n26306) );
  INVX1 U15244 ( .A(n29253), .Y(n26308) );
  INVX1 U15245 ( .A(n29253), .Y(n26309) );
  INVX1 U15246 ( .A(n29253), .Y(n26311) );
  INVX1 U15247 ( .A(n29253), .Y(n26312) );
  INVX1 U15248 ( .A(n29253), .Y(n26313) );
  INVX1 U15249 ( .A(n29253), .Y(n26315) );
  INVX1 U15250 ( .A(n29253), .Y(n26316) );
  INVX1 U15251 ( .A(n29253), .Y(n26317) );
  INVX1 U15252 ( .A(n29253), .Y(n26318) );
  INVX1 U15253 ( .A(n29253), .Y(n26319) );
  BUFX2 U15254 ( .A(n27276), .Y(n26320) );
  BUFX2 U15255 ( .A(n26306), .Y(n26321) );
  BUFX2 U15256 ( .A(n26306), .Y(n26322) );
  INVX1 U15257 ( .A(n26333), .Y(n26323) );
  INVX1 U15258 ( .A(n23202), .Y(n26325) );
  INVX1 U15259 ( .A(n26333), .Y(n26326) );
  INVX1 U15260 ( .A(n26332), .Y(n26328) );
  INVX1 U15261 ( .A(n26332), .Y(n26329) );
  INVX1 U15262 ( .A(n26325), .Y(n26330) );
  INVX1 U15263 ( .A(n26325), .Y(n26331) );
  INVX1 U15264 ( .A(n23202), .Y(n26332) );
  INVX1 U15265 ( .A(n23202), .Y(n26333) );
  INVX1 U15266 ( .A(n26332), .Y(n26334) );
  INVX1 U15267 ( .A(n26332), .Y(n26335) );
  INVX1 U15268 ( .A(n26333), .Y(n26336) );
  INVX1 U15269 ( .A(n34203), .Y(n26337) );
  INVX1 U15270 ( .A(n26337), .Y(n26338) );
  INVX1 U15271 ( .A(n28990), .Y(n26340) );
  BUFX2 U15272 ( .A(n28990), .Y(n26341) );
  BUFX2 U15273 ( .A(n28990), .Y(n26342) );
  INVX1 U15274 ( .A(n26341), .Y(n26343) );
  INVX1 U15275 ( .A(n26341), .Y(n26344) );
  INVX1 U15276 ( .A(n26341), .Y(n26345) );
  INVX1 U15277 ( .A(n26341), .Y(n26346) );
  INVX1 U15278 ( .A(n26341), .Y(n26347) );
  INVX1 U15279 ( .A(n26342), .Y(n26348) );
  INVX1 U15280 ( .A(n26342), .Y(n26349) );
  INVX1 U15281 ( .A(n26342), .Y(n26350) );
  INVX1 U15282 ( .A(n26342), .Y(n26351) );
  INVX1 U15283 ( .A(n26342), .Y(n26352) );
  BUFX2 U15284 ( .A(n28989), .Y(n26353) );
  BUFX2 U15285 ( .A(n28989), .Y(n26354) );
  INVX1 U15286 ( .A(n26353), .Y(n26355) );
  INVX1 U15287 ( .A(n26353), .Y(n26356) );
  INVX1 U15288 ( .A(n26353), .Y(n26357) );
  INVX1 U15289 ( .A(n26353), .Y(n26358) );
  INVX1 U15290 ( .A(n26353), .Y(n26359) );
  INVX1 U15291 ( .A(n26354), .Y(n26360) );
  INVX1 U15292 ( .A(n26354), .Y(n26361) );
  INVX1 U15293 ( .A(n26354), .Y(n26362) );
  INVX1 U15294 ( .A(n26354), .Y(n26363) );
  INVX1 U15295 ( .A(n26354), .Y(n26364) );
  BUFX2 U15296 ( .A(n29468), .Y(n26365) );
  BUFX2 U15297 ( .A(n29468), .Y(n26366) );
  INVX1 U15298 ( .A(n26365), .Y(n26367) );
  INVX1 U15299 ( .A(n26365), .Y(n26368) );
  INVX1 U15300 ( .A(n26365), .Y(n26369) );
  INVX1 U15301 ( .A(n26365), .Y(n26370) );
  INVX1 U15302 ( .A(n26365), .Y(n26371) );
  INVX1 U15303 ( .A(n26366), .Y(n26372) );
  INVX1 U15304 ( .A(n26366), .Y(n26373) );
  INVX1 U15305 ( .A(n26366), .Y(n26374) );
  INVX1 U15306 ( .A(n26366), .Y(n26375) );
  BUFX2 U15307 ( .A(n25703), .Y(n26376) );
  BUFX2 U15308 ( .A(n25703), .Y(n26377) );
  INVX1 U15309 ( .A(n26376), .Y(n26378) );
  INVX1 U15310 ( .A(n26376), .Y(n26379) );
  INVX1 U15311 ( .A(n26376), .Y(n26380) );
  INVX1 U15312 ( .A(n26376), .Y(n26381) );
  INVX1 U15313 ( .A(n26376), .Y(n26382) );
  INVX1 U15314 ( .A(n26377), .Y(n26383) );
  INVX1 U15315 ( .A(n26377), .Y(n26384) );
  INVX1 U15316 ( .A(n26377), .Y(n26385) );
  INVX1 U15317 ( .A(n26377), .Y(n26386) );
  INVX1 U15318 ( .A(n26377), .Y(n26387) );
  BUFX2 U15319 ( .A(n26366), .Y(n26388) );
  BUFX2 U15320 ( .A(n25703), .Y(n26389) );
  INVX1 U15321 ( .A(n26388), .Y(n26390) );
  INVX1 U15322 ( .A(n26388), .Y(n26391) );
  INVX1 U15323 ( .A(n26388), .Y(n26392) );
  INVX1 U15324 ( .A(n26388), .Y(n26393) );
  INVX1 U15325 ( .A(n26388), .Y(n26394) );
  INVX1 U15326 ( .A(n26389), .Y(n26395) );
  INVX1 U15327 ( .A(n26389), .Y(n26396) );
  INVX1 U15328 ( .A(n26389), .Y(n26397) );
  INVX1 U15329 ( .A(n26389), .Y(n26398) );
  INVX1 U15330 ( .A(n26389), .Y(n26399) );
  INVX1 U15331 ( .A(n25704), .Y(n26400) );
  INVX1 U15332 ( .A(n25704), .Y(n26401) );
  INVX1 U15333 ( .A(n25704), .Y(n26402) );
  INVX1 U15334 ( .A(n25704), .Y(n26403) );
  INVX1 U15335 ( .A(n25704), .Y(n26404) );
  INVX1 U15336 ( .A(n26400), .Y(n26405) );
  INVX1 U15337 ( .A(n26400), .Y(n26406) );
  INVX1 U15338 ( .A(n26400), .Y(n26407) );
  INVX1 U15339 ( .A(n26400), .Y(n26408) );
  INVX1 U15340 ( .A(n26401), .Y(n26409) );
  INVX1 U15341 ( .A(n26401), .Y(n26410) );
  INVX1 U15342 ( .A(n26401), .Y(n26411) );
  INVX1 U15343 ( .A(n26402), .Y(n26412) );
  INVX1 U15344 ( .A(n26402), .Y(n26413) );
  INVX1 U15345 ( .A(n26402), .Y(n26414) );
  INVX1 U15346 ( .A(n26402), .Y(n26415) );
  INVX1 U15347 ( .A(n26403), .Y(n26416) );
  INVX1 U15348 ( .A(n26403), .Y(n26417) );
  INVX1 U15349 ( .A(n26403), .Y(n26418) );
  INVX1 U15350 ( .A(n26403), .Y(n26419) );
  INVX1 U15351 ( .A(n26404), .Y(n26420) );
  INVX1 U15352 ( .A(n26404), .Y(n26421) );
  INVX1 U15353 ( .A(n26404), .Y(n26422) );
  INVX1 U15354 ( .A(n26340), .Y(n26423) );
  INVX1 U15355 ( .A(n26340), .Y(n26424) );
  INVX1 U15356 ( .A(n26340), .Y(n26425) );
  INVX1 U15357 ( .A(n26340), .Y(n26426) );
  INVX1 U15358 ( .A(n26423), .Y(n26427) );
  INVX1 U15359 ( .A(n26423), .Y(n26428) );
  INVX1 U15360 ( .A(n26423), .Y(n26429) );
  INVX1 U15361 ( .A(n26423), .Y(n26430) );
  INVX1 U15362 ( .A(n26424), .Y(n26431) );
  INVX1 U15363 ( .A(n26424), .Y(n26432) );
  INVX1 U15364 ( .A(n26424), .Y(n26433) );
  INVX1 U15365 ( .A(n26424), .Y(n26434) );
  INVX1 U15366 ( .A(n26425), .Y(n26435) );
  INVX1 U15367 ( .A(n26425), .Y(n26436) );
  INVX1 U15368 ( .A(n26425), .Y(n26437) );
  INVX1 U15369 ( .A(n26425), .Y(n26438) );
  INVX1 U15370 ( .A(n26426), .Y(n26439) );
  INVX1 U15371 ( .A(n26426), .Y(n26440) );
  INVX1 U15372 ( .A(n26426), .Y(n26441) );
  INVX1 U15373 ( .A(n26426), .Y(n26442) );
  INVX1 U15374 ( .A(n26365), .Y(n26443) );
  INVX1 U15375 ( .A(n26404), .Y(n26444) );
  INVX2 U15376 ( .A(n2246), .Y(n29468) );
  INVX1 U15377 ( .A(n26450), .Y(n26447) );
  INVX1 U15378 ( .A(n29231), .Y(n26448) );
  INVX1 U15379 ( .A(n26464), .Y(n26449) );
  BUFX2 U15380 ( .A(n26463), .Y(n26450) );
  BUFX2 U15381 ( .A(n29231), .Y(n26451) );
  BUFX2 U15382 ( .A(n26463), .Y(n26452) );
  INVX1 U15383 ( .A(n26450), .Y(n26453) );
  INVX1 U15384 ( .A(n26450), .Y(n26454) );
  INVX1 U15385 ( .A(n26451), .Y(n26455) );
  INVX1 U15386 ( .A(n26451), .Y(n26456) );
  INVX1 U15387 ( .A(n26451), .Y(n26457) );
  INVX1 U15388 ( .A(n26451), .Y(n26458) );
  INVX1 U15389 ( .A(n26452), .Y(n26459) );
  INVX1 U15390 ( .A(n26452), .Y(n26460) );
  INVX1 U15391 ( .A(n26452), .Y(n26461) );
  INVX1 U15392 ( .A(n26452), .Y(n26462) );
  INVX1 U15393 ( .A(n26464), .Y(n26465) );
  INVX1 U15394 ( .A(n26464), .Y(n26466) );
  INVX1 U15395 ( .A(n26464), .Y(n26467) );
  INVX1 U15396 ( .A(n26463), .Y(n26468) );
  INVX1 U15397 ( .A(n26464), .Y(n26469) );
  INVX1 U15398 ( .A(n26463), .Y(n26470) );
  INVX1 U15399 ( .A(n26464), .Y(n26471) );
  INVX1 U15400 ( .A(n26463), .Y(n26472) );
  INVX1 U15401 ( .A(n26464), .Y(n26473) );
  INVX1 U15402 ( .A(n26463), .Y(n26474) );
  INVX1 U15403 ( .A(n26463), .Y(n26475) );
  INVX1 U15404 ( .A(n26463), .Y(n26476) );
  INVX1 U15405 ( .A(n26464), .Y(n26477) );
  INVX1 U15406 ( .A(n29231), .Y(n26478) );
  INVX1 U15407 ( .A(n26464), .Y(n26479) );
  AND2X2 U15408 ( .A(n30637), .B(n30636), .Y(n27299) );
  AND2X2 U15409 ( .A(n23295), .B(n29331), .Y(n27220) );
  INVX1 U15410 ( .A(n2250), .Y(n26480) );
  INVX1 U15411 ( .A(n26480), .Y(n26481) );
  INVX1 U15412 ( .A(n26480), .Y(n26482) );
  AND2X2 U15413 ( .A(n23293), .B(n29331), .Y(n27219) );
  INVX4 U15414 ( .A(n26941), .Y(n33718) );
  INVX8 U15415 ( .A(n26878), .Y(n34222) );
  INVX2 U15416 ( .A(n34218), .Y(n26878) );
  INVX8 U15417 ( .A(n23611), .Y(n29683) );
  AND2X2 U15418 ( .A(n23440), .B(n23611), .Y(n27301) );
  AND2X2 U15419 ( .A(n23289), .B(n29331), .Y(n27225) );
  INVX4 U15420 ( .A(n27253), .Y(n29330) );
  INVX1 U15421 ( .A(n21073), .Y(n26485) );
  INVX1 U15422 ( .A(n21095), .Y(n26486) );
  INVX1 U15423 ( .A(n21095), .Y(n26487) );
  INVX1 U15424 ( .A(n21095), .Y(n26488) );
  INVX1 U15425 ( .A(n21095), .Y(n26489) );
  INVX1 U15426 ( .A(n21095), .Y(n26490) );
  INVX1 U15427 ( .A(n21095), .Y(n26491) );
  INVX1 U15428 ( .A(n21095), .Y(n26492) );
  INVX1 U15429 ( .A(n28599), .Y(n26493) );
  INVX1 U15430 ( .A(n28599), .Y(n26494) );
  INVX1 U15431 ( .A(n28599), .Y(n26495) );
  INVX1 U15432 ( .A(n28599), .Y(n26496) );
  INVX1 U15433 ( .A(n28599), .Y(n26497) );
  INVX1 U15434 ( .A(n28599), .Y(n26498) );
  INVX1 U15435 ( .A(n28599), .Y(n26499) );
  INVX1 U15436 ( .A(n26514), .Y(n26501) );
  INVX1 U15437 ( .A(n26514), .Y(n26502) );
  INVX1 U15438 ( .A(n26514), .Y(n26503) );
  INVX1 U15439 ( .A(n28600), .Y(n26505) );
  INVX1 U15440 ( .A(n28600), .Y(n26506) );
  INVX1 U15441 ( .A(n28600), .Y(n26507) );
  INVX1 U15442 ( .A(n28600), .Y(n26508) );
  INVX1 U15443 ( .A(n21073), .Y(n26509) );
  INVX1 U15444 ( .A(n28601), .Y(n26510) );
  INVX1 U15445 ( .A(n28601), .Y(n26511) );
  INVX1 U15446 ( .A(n21073), .Y(n26512) );
  INVX1 U15447 ( .A(n21073), .Y(n26513) );
  AND2X2 U15448 ( .A(n29807), .B(n25724), .Y(n27218) );
  INVX4 U15449 ( .A(n23109), .Y(n32491) );
  INVX4 U15450 ( .A(n27194), .Y(n33216) );
  INVX1 U15451 ( .A(net89777), .Y(net106017) );
  INVX1 U15452 ( .A(net106017), .Y(net106018) );
  INVX4 U15453 ( .A(n22947), .Y(n26518) );
  BUFX4 U15454 ( .A(n25743), .Y(n26519) );
  INVX1 U15455 ( .A(n26078), .Y(n26520) );
  INVX1 U15456 ( .A(n28991), .Y(n26522) );
  BUFX2 U15457 ( .A(n28991), .Y(n26523) );
  BUFX2 U15458 ( .A(n28991), .Y(n26524) );
  INVX1 U15459 ( .A(n26523), .Y(n26525) );
  INVX1 U15460 ( .A(n26523), .Y(n26526) );
  INVX1 U15461 ( .A(n26523), .Y(n26527) );
  INVX1 U15462 ( .A(n26523), .Y(n26528) );
  INVX1 U15463 ( .A(n26523), .Y(n26529) );
  INVX1 U15464 ( .A(n26524), .Y(n26530) );
  INVX1 U15465 ( .A(n26524), .Y(n26531) );
  INVX1 U15466 ( .A(n26524), .Y(n26532) );
  INVX1 U15467 ( .A(n26524), .Y(n26533) );
  INVX1 U15468 ( .A(n26524), .Y(n26534) );
  BUFX2 U15469 ( .A(n29466), .Y(n26535) );
  BUFX2 U15470 ( .A(n29466), .Y(n26536) );
  INVX1 U15471 ( .A(n26535), .Y(n26537) );
  INVX1 U15472 ( .A(n26535), .Y(n26538) );
  INVX1 U15473 ( .A(n26535), .Y(n26539) );
  INVX1 U15474 ( .A(n26535), .Y(n26540) );
  INVX1 U15475 ( .A(n26535), .Y(n26541) );
  INVX1 U15476 ( .A(n26536), .Y(n26542) );
  INVX1 U15477 ( .A(n26536), .Y(n26543) );
  INVX1 U15478 ( .A(n26536), .Y(n26544) );
  INVX1 U15479 ( .A(n26536), .Y(n26545) );
  INVX1 U15480 ( .A(n26536), .Y(n26546) );
  BUFX2 U15481 ( .A(n26047), .Y(n26547) );
  BUFX2 U15482 ( .A(n26047), .Y(n26548) );
  INVX1 U15483 ( .A(n26547), .Y(n26549) );
  INVX1 U15484 ( .A(n26547), .Y(n26550) );
  INVX1 U15485 ( .A(n26547), .Y(n26551) );
  INVX1 U15486 ( .A(n26547), .Y(n26552) );
  INVX1 U15487 ( .A(n26547), .Y(n26553) );
  INVX1 U15488 ( .A(n26548), .Y(n26554) );
  INVX1 U15489 ( .A(n26548), .Y(n26555) );
  INVX1 U15490 ( .A(n26548), .Y(n26556) );
  INVX1 U15491 ( .A(n26548), .Y(n26557) );
  INVX1 U15492 ( .A(n26548), .Y(n26558) );
  INVX1 U15493 ( .A(n26048), .Y(n26559) );
  INVX1 U15494 ( .A(n26048), .Y(n26560) );
  INVX1 U15495 ( .A(n26048), .Y(n26561) );
  INVX1 U15496 ( .A(n26559), .Y(n26562) );
  INVX1 U15497 ( .A(n26559), .Y(n26563) );
  INVX1 U15498 ( .A(n26559), .Y(n26564) );
  INVX1 U15499 ( .A(n26560), .Y(n26565) );
  INVX1 U15500 ( .A(n26560), .Y(n26566) );
  INVX1 U15501 ( .A(n26560), .Y(n26567) );
  INVX1 U15502 ( .A(n26560), .Y(n26568) );
  INVX1 U15503 ( .A(n26561), .Y(n26569) );
  INVX1 U15504 ( .A(n26561), .Y(n26570) );
  INVX1 U15505 ( .A(n26561), .Y(n26571) );
  INVX1 U15506 ( .A(n26561), .Y(n26572) );
  INVX1 U15507 ( .A(n26522), .Y(n26573) );
  INVX1 U15508 ( .A(n26573), .Y(n26574) );
  INVX1 U15509 ( .A(n26573), .Y(n26575) );
  INVX1 U15510 ( .A(n26573), .Y(n26576) );
  INVX8 U15511 ( .A(n27175), .Y(n30626) );
  INVX8 U15512 ( .A(net105857), .Y(net105859) );
  INVX1 U15513 ( .A(net113687), .Y(net105793) );
  INVX1 U15514 ( .A(net113687), .Y(net105794) );
  INVX1 U15515 ( .A(net149877), .Y(net105797) );
  INVX1 U15516 ( .A(net149876), .Y(net105801) );
  INVX1 U15517 ( .A(net113687), .Y(net105802) );
  INVX1 U15518 ( .A(alt14_net96326), .Y(net105808) );
  INVX1 U15519 ( .A(net149877), .Y(net105816) );
  OR2X1 U15520 ( .A(n29368), .B(n34132), .Y(n21742) );
  INVX1 U15521 ( .A(n21742), .Y(n26577) );
  OR2X1 U15522 ( .A(n29367), .B(n34119), .Y(n21729) );
  INVX1 U15523 ( .A(n21729), .Y(n26578) );
  OR2X1 U15524 ( .A(n29366), .B(n34106), .Y(n21716) );
  INVX1 U15525 ( .A(n21716), .Y(n26579) );
  OR2X1 U15526 ( .A(n29370), .B(n34158), .Y(n21769) );
  INVX1 U15527 ( .A(n21769), .Y(n26580) );
  INVX1 U15528 ( .A(n21755), .Y(n26581) );
  OR2X1 U15529 ( .A(n29371), .B(n34093), .Y(n21703) );
  INVX1 U15530 ( .A(n21703), .Y(n26582) );
  OR2X1 U15531 ( .A(n29371), .B(n34080), .Y(n21689) );
  INVX1 U15532 ( .A(n21689), .Y(n26583) );
  OR2X1 U15533 ( .A(n29370), .B(n34067), .Y(n21676) );
  INVX1 U15534 ( .A(n21676), .Y(n26584) );
  OR2X1 U15535 ( .A(n29365), .B(n34054), .Y(n21662) );
  INVX1 U15536 ( .A(n21662), .Y(n26585) );
  OR2X1 U15537 ( .A(n29370), .B(n34041), .Y(n21649) );
  INVX1 U15538 ( .A(n21649), .Y(n26586) );
  OR2X1 U15539 ( .A(n29370), .B(n34028), .Y(n21636) );
  INVX1 U15540 ( .A(n21636), .Y(n26587) );
  BUFX2 U15541 ( .A(n14396), .Y(n26588) );
  BUFX2 U15542 ( .A(n14489), .Y(n26589) );
  BUFX2 U15543 ( .A(n14659), .Y(n26590) );
  BUFX2 U15544 ( .A(n14832), .Y(n26591) );
  BUFX2 U15545 ( .A(n15004), .Y(n26592) );
  AND2X1 U15546 ( .A(n29221), .B(n27170), .Y(n30655) );
  INVX1 U15547 ( .A(n30655), .Y(n26593) );
  AND2X1 U15548 ( .A(n27273), .B(n29775), .Y(n30500) );
  INVX1 U15549 ( .A(n30500), .Y(n26594) );
  INVX1 U15550 ( .A(n31882), .Y(n26595) );
  INVX1 U15551 ( .A(n31511), .Y(n26596) );
  INVX1 U15552 ( .A(n31259), .Y(n26597) );
  OR2X1 U15553 ( .A(n29371), .B(n34229), .Y(n21781) );
  INVX1 U15554 ( .A(n21781), .Y(n26598) );
  OR2X1 U15555 ( .A(n29368), .B(n34131), .Y(n21741) );
  INVX1 U15556 ( .A(n21741), .Y(n26599) );
  OR2X1 U15557 ( .A(n29367), .B(n34118), .Y(n21728) );
  INVX1 U15558 ( .A(n21728), .Y(n26600) );
  OR2X1 U15559 ( .A(n29366), .B(n34105), .Y(n21715) );
  INVX1 U15560 ( .A(n21715), .Y(n26601) );
  OR2X1 U15561 ( .A(n29370), .B(n34157), .Y(n21768) );
  INVX1 U15562 ( .A(n21768), .Y(n26602) );
  INVX1 U15563 ( .A(n21754), .Y(n26603) );
  OR2X1 U15564 ( .A(n29371), .B(n34092), .Y(n21702) );
  INVX1 U15565 ( .A(n21702), .Y(n26604) );
  OR2X1 U15566 ( .A(n29371), .B(n34079), .Y(n21688) );
  INVX1 U15567 ( .A(n21688), .Y(n26605) );
  OR2X1 U15568 ( .A(n29370), .B(n34066), .Y(n21675) );
  INVX1 U15569 ( .A(n21675), .Y(n26606) );
  OR2X1 U15570 ( .A(n29365), .B(n34053), .Y(n21661) );
  INVX1 U15571 ( .A(n21661), .Y(n26607) );
  OR2X1 U15572 ( .A(n29370), .B(n34040), .Y(n21648) );
  INVX1 U15573 ( .A(n21648), .Y(n26608) );
  OR2X1 U15574 ( .A(n29370), .B(n34027), .Y(n21635) );
  INVX1 U15575 ( .A(n21635), .Y(n26609) );
  OR2X2 U15576 ( .A(n21089), .B(n29363), .Y(n21599) );
  INVX1 U15577 ( .A(n21599), .Y(n26610) );
  OR2X1 U15578 ( .A(n29364), .B(n34016), .Y(n21624) );
  INVX1 U15579 ( .A(n21624), .Y(n26611) );
  AND2X1 U15580 ( .A(n16236), .B(n16233), .Y(n16235) );
  INVX1 U15581 ( .A(n16235), .Y(n26612) );
  BUFX2 U15582 ( .A(n14422), .Y(n26613) );
  BUFX2 U15583 ( .A(n14513), .Y(n26614) );
  BUFX2 U15584 ( .A(n14671), .Y(n26615) );
  BUFX2 U15585 ( .A(n14856), .Y(n26616) );
  BUFX2 U15586 ( .A(n15028), .Y(n26617) );
  AND2X2 U15587 ( .A(n29352), .B(n30508), .Y(n29790) );
  INVX1 U15588 ( .A(n29790), .Y(n26618) );
  AND2X1 U15589 ( .A(n27273), .B(n29783), .Y(n30505) );
  INVX1 U15590 ( .A(n30505), .Y(n26619) );
  INVX1 U15591 ( .A(n31841), .Y(n26620) );
  AND2X1 U15592 ( .A(n29221), .B(n26926), .Y(n31492) );
  INVX1 U15593 ( .A(n31492), .Y(n26621) );
  INVX1 U15594 ( .A(n31219), .Y(n26622) );
  INVX1 U15595 ( .A(n30886), .Y(n26623) );
  OR2X1 U15596 ( .A(n29371), .B(n34169), .Y(n21780) );
  INVX1 U15597 ( .A(n21780), .Y(n26624) );
  OR2X1 U15598 ( .A(n29368), .B(n34130), .Y(n21740) );
  INVX1 U15599 ( .A(n21740), .Y(n26625) );
  OR2X1 U15600 ( .A(n29367), .B(n34117), .Y(n21727) );
  INVX1 U15601 ( .A(n21727), .Y(n26626) );
  OR2X1 U15602 ( .A(n29366), .B(n34104), .Y(n21714) );
  INVX1 U15603 ( .A(n21714), .Y(n26627) );
  OR2X1 U15604 ( .A(n29370), .B(n34156), .Y(n21766) );
  INVX1 U15605 ( .A(n21766), .Y(n26628) );
  INVX1 U15606 ( .A(n21753), .Y(n26629) );
  OR2X1 U15607 ( .A(n29371), .B(n34091), .Y(n21701) );
  INVX1 U15608 ( .A(n21701), .Y(n26630) );
  OR2X1 U15609 ( .A(n29371), .B(n34078), .Y(n21687) );
  INVX1 U15610 ( .A(n21687), .Y(n26631) );
  OR2X1 U15611 ( .A(n29370), .B(n34065), .Y(n21674) );
  INVX1 U15612 ( .A(n21674), .Y(n26632) );
  OR2X1 U15613 ( .A(n29365), .B(n34052), .Y(n21660) );
  INVX1 U15614 ( .A(n21660), .Y(n26633) );
  OR2X1 U15615 ( .A(n29370), .B(n34039), .Y(n21647) );
  INVX1 U15616 ( .A(n21647), .Y(n26634) );
  OR2X1 U15617 ( .A(n29370), .B(n34026), .Y(n21634) );
  INVX1 U15618 ( .A(n21634), .Y(n26635) );
  OR2X2 U15619 ( .A(n29461), .B(n29363), .Y(n21602) );
  INVX1 U15620 ( .A(n21602), .Y(n26636) );
  OR2X1 U15621 ( .A(n29364), .B(n34015), .Y(n21623) );
  INVX1 U15622 ( .A(n21623), .Y(n26637) );
  AND2X1 U15623 ( .A(n16245), .B(n16242), .Y(n16244) );
  INVX1 U15624 ( .A(n16244), .Y(n26638) );
  BUFX2 U15625 ( .A(n14435), .Y(n26639) );
  BUFX2 U15626 ( .A(n14501), .Y(n26640) );
  BUFX2 U15627 ( .A(n14710), .Y(n26641) );
  BUFX2 U15628 ( .A(n14868), .Y(n26642) );
  BUFX2 U15629 ( .A(n15040), .Y(n26643) );
  AND2X2 U15630 ( .A(n29352), .B(n30513), .Y(n29799) );
  INVX1 U15631 ( .A(n29799), .Y(n26644) );
  AND2X1 U15632 ( .A(n27273), .B(n29791), .Y(n30510) );
  INVX1 U15633 ( .A(n30510), .Y(n26645) );
  INVX1 U15634 ( .A(n31802), .Y(n26646) );
  INVX1 U15635 ( .A(n31473), .Y(n26647) );
  INVX1 U15636 ( .A(n31179), .Y(n26648) );
  AND2X1 U15637 ( .A(n29221), .B(n27169), .Y(n30865) );
  INVX1 U15638 ( .A(n30865), .Y(n26649) );
  OR2X1 U15639 ( .A(n29371), .B(n34168), .Y(n21779) );
  INVX1 U15640 ( .A(n21779), .Y(n26650) );
  OR2X1 U15641 ( .A(n29368), .B(n34129), .Y(n21739) );
  INVX1 U15642 ( .A(n21739), .Y(n26651) );
  OR2X1 U15643 ( .A(n29367), .B(n34116), .Y(n21726) );
  INVX1 U15644 ( .A(n21726), .Y(n26652) );
  OR2X1 U15645 ( .A(n29366), .B(n34103), .Y(n21713) );
  INVX1 U15646 ( .A(n21713), .Y(n26653) );
  OR2X1 U15647 ( .A(n29370), .B(n34155), .Y(n21765) );
  INVX1 U15648 ( .A(n21765), .Y(n26654) );
  INVX1 U15649 ( .A(n21752), .Y(n26655) );
  OR2X1 U15650 ( .A(n29371), .B(n34090), .Y(n21700) );
  INVX1 U15651 ( .A(n21700), .Y(n26656) );
  OR2X1 U15652 ( .A(n29371), .B(n34077), .Y(n21686) );
  INVX1 U15653 ( .A(n21686), .Y(n26657) );
  OR2X1 U15654 ( .A(n29370), .B(n34064), .Y(n21673) );
  INVX1 U15655 ( .A(n21673), .Y(n26658) );
  OR2X1 U15656 ( .A(n29365), .B(n34051), .Y(n21659) );
  INVX1 U15657 ( .A(n21659), .Y(n26659) );
  OR2X1 U15658 ( .A(n29370), .B(n34038), .Y(n21646) );
  INVX1 U15659 ( .A(n21646), .Y(n26660) );
  OR2X1 U15660 ( .A(n29370), .B(n34025), .Y(n21633) );
  INVX1 U15661 ( .A(n21633), .Y(n26661) );
  OR2X2 U15662 ( .A(n26515), .B(n29363), .Y(n21600) );
  INVX1 U15663 ( .A(n21600), .Y(n26662) );
  OR2X1 U15664 ( .A(n29364), .B(n34014), .Y(n21622) );
  INVX1 U15665 ( .A(n21622), .Y(n26663) );
  AND2X1 U15666 ( .A(n29640), .B(n29639), .Y(n29641) );
  INVX1 U15667 ( .A(n29641), .Y(n26664) );
  BUFX2 U15668 ( .A(n16153), .Y(n26665) );
  BUFX2 U15669 ( .A(n16155), .Y(n26666) );
  OR2X2 U15670 ( .A(nc[19]), .B(nc[18]), .Y(n29532) );
  INVX1 U15671 ( .A(n29532), .Y(n26667) );
  BUFX2 U15672 ( .A(n29636), .Y(n26668) );
  BUFX2 U15673 ( .A(n14537), .Y(n26669) );
  BUFX2 U15674 ( .A(n14722), .Y(n26670) );
  BUFX2 U15675 ( .A(n14894), .Y(n26671) );
  BUFX2 U15676 ( .A(n15052), .Y(n26672) );
  BUFX2 U15677 ( .A(n15077), .Y(n26673) );
  AND2X1 U15678 ( .A(n30319), .B(n30457), .Y(n31380) );
  INVX1 U15679 ( .A(n31380), .Y(n26674) );
  AND2X1 U15680 ( .A(n30135), .B(n27323), .Y(n30793) );
  INVX1 U15681 ( .A(n30793), .Y(n26675) );
  AND2X2 U15682 ( .A(n29352), .B(n30531), .Y(n29841) );
  INVX1 U15683 ( .A(n29841), .Y(n26676) );
  AND2X1 U15684 ( .A(n27273), .B(n29800), .Y(n30515) );
  INVX1 U15685 ( .A(n30515), .Y(n26677) );
  INVX1 U15686 ( .A(n31762), .Y(n26678) );
  AND2X1 U15687 ( .A(n29221), .B(n26991), .Y(n31453) );
  INVX1 U15688 ( .A(n31453), .Y(n26679) );
  INVX1 U15689 ( .A(n31142), .Y(n26680) );
  INVX1 U15690 ( .A(n30846), .Y(n26681) );
  OR2X1 U15691 ( .A(n29371), .B(n34167), .Y(n21778) );
  INVX1 U15692 ( .A(n21778), .Y(n26682) );
  OR2X1 U15693 ( .A(n29368), .B(n34128), .Y(n21738) );
  INVX1 U15694 ( .A(n21738), .Y(n26683) );
  OR2X1 U15695 ( .A(n29367), .B(n34115), .Y(n21725) );
  INVX1 U15696 ( .A(n21725), .Y(n26684) );
  OR2X1 U15697 ( .A(n29366), .B(n34102), .Y(n21712) );
  INVX1 U15698 ( .A(n21712), .Y(n26685) );
  OR2X1 U15699 ( .A(n29370), .B(n34154), .Y(n21764) );
  INVX1 U15700 ( .A(n21764), .Y(n26686) );
  INVX1 U15701 ( .A(n21751), .Y(n26687) );
  OR2X1 U15702 ( .A(n29371), .B(n34089), .Y(n21698) );
  INVX1 U15703 ( .A(n21698), .Y(n26688) );
  OR2X1 U15704 ( .A(n29371), .B(n34076), .Y(n21685) );
  INVX1 U15705 ( .A(n21685), .Y(n26689) );
  OR2X1 U15706 ( .A(n29370), .B(n34063), .Y(n21672) );
  INVX1 U15707 ( .A(n21672), .Y(n26690) );
  OR2X1 U15708 ( .A(n29365), .B(n34050), .Y(n21658) );
  INVX1 U15709 ( .A(n21658), .Y(n26691) );
  OR2X1 U15710 ( .A(n29371), .B(n34037), .Y(n21645) );
  INVX1 U15711 ( .A(n21645), .Y(n26692) );
  OR2X1 U15712 ( .A(n29370), .B(n34024), .Y(n21632) );
  INVX1 U15713 ( .A(n21632), .Y(n26693) );
  OR2X2 U15714 ( .A(n28603), .B(n29363), .Y(n21601) );
  INVX1 U15715 ( .A(n21601), .Y(n26694) );
  OR2X1 U15716 ( .A(n29364), .B(n34013), .Y(n21621) );
  INVX1 U15717 ( .A(n21621), .Y(n26695) );
  AND2X1 U15718 ( .A(n16032), .B(n34567), .Y(n16031) );
  INVX1 U15719 ( .A(n16031), .Y(n26696) );
  OR2X2 U15720 ( .A(nc[4]), .B(nc[3]), .Y(n29549) );
  INVX1 U15721 ( .A(n29549), .Y(n26697) );
  AND2X1 U15722 ( .A(n27274), .B(n16242), .Y(n16229) );
  INVX1 U15723 ( .A(n16229), .Y(n26698) );
  BUFX2 U15724 ( .A(n16230), .Y(n26699) );
  OR2X1 U15725 ( .A(n27007), .B(n27184), .Y(n16231) );
  BUFX2 U15726 ( .A(n14474), .Y(n26700) );
  BUFX2 U15727 ( .A(n14525), .Y(n26701) );
  BUFX2 U15728 ( .A(n14734), .Y(n26702) );
  BUFX2 U15729 ( .A(n14906), .Y(n26703) );
  BUFX2 U15730 ( .A(n15089), .Y(n26704) );
  AND2X1 U15731 ( .A(n30409), .B(n30432), .Y(n31635) );
  INVX1 U15732 ( .A(n31635), .Y(n26705) );
  AND2X1 U15733 ( .A(n30135), .B(n30457), .Y(n30753) );
  INVX1 U15734 ( .A(n30753), .Y(n26706) );
  AND2X2 U15735 ( .A(n29352), .B(n30535), .Y(n29851) );
  INVX1 U15736 ( .A(n29851), .Y(n26707) );
  AND2X1 U15737 ( .A(n30038), .B(n29730), .Y(n29750) );
  INVX1 U15738 ( .A(n29750), .Y(n26708) );
  AND2X1 U15739 ( .A(n27273), .B(n29812), .Y(n30520) );
  INVX1 U15740 ( .A(n30520), .Y(n26709) );
  AND2X2 U15741 ( .A(n29831), .B(n27314), .Y(n29933) );
  INVX1 U15742 ( .A(n29933), .Y(n26710) );
  INVX1 U15743 ( .A(n31724), .Y(n26711) );
  INVX1 U15744 ( .A(n31434), .Y(n26712) );
  INVX1 U15745 ( .A(n31102), .Y(n26713) );
  AND2X1 U15746 ( .A(n29221), .B(n27072), .Y(n30825) );
  INVX1 U15747 ( .A(n30825), .Y(n26714) );
  AND2X2 U15748 ( .A(n27236), .B(n27239), .Y(n31959) );
  INVX1 U15749 ( .A(n31959), .Y(n26715) );
  INVX1 U15750 ( .A(n31959), .Y(n26716) );
  OR2X1 U15751 ( .A(n29371), .B(n34166), .Y(n21777) );
  INVX1 U15752 ( .A(n21777), .Y(n26717) );
  OR2X1 U15753 ( .A(n29368), .B(n34127), .Y(n21737) );
  INVX1 U15754 ( .A(n21737), .Y(n26718) );
  OR2X1 U15755 ( .A(n29367), .B(n34114), .Y(n21724) );
  INVX1 U15756 ( .A(n21724), .Y(n26719) );
  OR2X1 U15757 ( .A(n29366), .B(n34101), .Y(n21711) );
  INVX1 U15758 ( .A(n21711), .Y(n26720) );
  OR2X1 U15759 ( .A(n29370), .B(n34153), .Y(n21763) );
  INVX1 U15760 ( .A(n21763), .Y(n26721) );
  INVX1 U15761 ( .A(n21750), .Y(n26722) );
  OR2X1 U15762 ( .A(n29371), .B(n34088), .Y(n21697) );
  INVX1 U15763 ( .A(n21697), .Y(n26723) );
  OR2X1 U15764 ( .A(n29371), .B(n34075), .Y(n21684) );
  INVX1 U15765 ( .A(n21684), .Y(n26724) );
  OR2X1 U15766 ( .A(n29370), .B(n34062), .Y(n21671) );
  INVX1 U15767 ( .A(n21671), .Y(n26725) );
  OR2X1 U15768 ( .A(n29365), .B(n34049), .Y(n21657) );
  INVX1 U15769 ( .A(n21657), .Y(n26726) );
  OR2X1 U15770 ( .A(n29370), .B(n34036), .Y(n21644) );
  INVX1 U15771 ( .A(n21644), .Y(n26727) );
  OR2X1 U15772 ( .A(n29370), .B(n34023), .Y(n21631) );
  INVX1 U15773 ( .A(n21631), .Y(n26728) );
  OR2X2 U15774 ( .A(n33996), .B(n29363), .Y(n21604) );
  INVX1 U15775 ( .A(n21604), .Y(n26729) );
  OR2X1 U15776 ( .A(n29364), .B(n34012), .Y(n21620) );
  INVX1 U15777 ( .A(n21620), .Y(n26730) );
  AND2X1 U15778 ( .A(n16190), .B(n34561), .Y(n16189) );
  INVX1 U15779 ( .A(n16189), .Y(n26731) );
  BUFX2 U15780 ( .A(n16002), .Y(n26732) );
  BUFX2 U15781 ( .A(n16004), .Y(n26733) );
  AND2X1 U15782 ( .A(n16224), .B(n29654), .Y(n16217) );
  INVX1 U15783 ( .A(n16217), .Y(n26734) );
  BUFX2 U15784 ( .A(n29736), .Y(n26735) );
  BUFX2 U15785 ( .A(n29546), .Y(n26736) );
  OR2X2 U15786 ( .A(nc[12]), .B(nc[11]), .Y(n29543) );
  INVX1 U15787 ( .A(n29543), .Y(n26737) );
  BUFX2 U15788 ( .A(n14461), .Y(n26738) );
  BUFX2 U15789 ( .A(n14573), .Y(n26739) );
  BUFX2 U15790 ( .A(n14746), .Y(n26740) );
  BUFX2 U15791 ( .A(n14918), .Y(n26741) );
  BUFX2 U15792 ( .A(n15101), .Y(n26742) );
  AND2X1 U15793 ( .A(n30409), .B(n30418), .Y(n31598) );
  INVX1 U15794 ( .A(n31598), .Y(n26743) );
  AND2X1 U15795 ( .A(n30319), .B(n30426), .Y(n31303) );
  INVX1 U15796 ( .A(n31303), .Y(n26744) );
  AND2X1 U15797 ( .A(n30225), .B(n30432), .Y(n31011) );
  INVX1 U15798 ( .A(n31011), .Y(n26745) );
  AND2X1 U15799 ( .A(n30135), .B(n30440), .Y(n30713) );
  INVX1 U15800 ( .A(n30713), .Y(n26746) );
  AND2X2 U15801 ( .A(n29352), .B(n30489), .Y(n29754) );
  INVX1 U15802 ( .A(n29754), .Y(n26747) );
  AND2X2 U15803 ( .A(n29352), .B(n30545), .Y(n29867) );
  INVX1 U15804 ( .A(n29867), .Y(n26748) );
  AND2X1 U15805 ( .A(n27274), .B(n26859), .Y(n16015) );
  INVX1 U15806 ( .A(n16015), .Y(n26749) );
  AND2X2 U15807 ( .A(n29352), .B(n30586), .Y(n29961) );
  INVX1 U15808 ( .A(n29961), .Y(n26750) );
  AND2X1 U15809 ( .A(n27273), .B(n29832), .Y(n30528) );
  INVX1 U15810 ( .A(n30528), .Y(n26751) );
  AND2X2 U15811 ( .A(n30012), .B(n27314), .Y(n29922) );
  INVX1 U15812 ( .A(n29922), .Y(n26752) );
  AND2X2 U15813 ( .A(n30281), .B(T[4]), .Y(n29644) );
  INVX1 U15814 ( .A(n29644), .Y(n26753) );
  INVX4 U15815 ( .A(n26272), .Y(n30281) );
  INVX1 U15816 ( .A(n31685), .Y(n26754) );
  AND2X1 U15817 ( .A(n29221), .B(n26927), .Y(n31413) );
  INVX1 U15818 ( .A(n31413), .Y(n26755) );
  INVX1 U15819 ( .A(n31062), .Y(n26756) );
  INVX1 U15820 ( .A(n30806), .Y(n26757) );
  AND2X2 U15821 ( .A(n30227), .B(n30442), .Y(n32005) );
  INVX1 U15822 ( .A(n32005), .Y(n26758) );
  INVX1 U15823 ( .A(n32005), .Y(n26759) );
  AND2X2 U15824 ( .A(n27265), .B(n30458), .Y(n31943) );
  INVX1 U15825 ( .A(n31943), .Y(n26760) );
  INVX1 U15826 ( .A(n31943), .Y(n26761) );
  AND2X2 U15827 ( .A(n27236), .B(n27237), .Y(n31964) );
  INVX1 U15828 ( .A(n31964), .Y(n26762) );
  INVX1 U15829 ( .A(n31964), .Y(n26763) );
  AND2X2 U15830 ( .A(n29835), .B(n30040), .Y(n33726) );
  INVX1 U15831 ( .A(n33726), .Y(n26765) );
  OR2X1 U15832 ( .A(n29371), .B(n34165), .Y(n21776) );
  INVX1 U15833 ( .A(n21776), .Y(n26766) );
  OR2X1 U15834 ( .A(n29368), .B(n34126), .Y(n21736) );
  INVX1 U15835 ( .A(n21736), .Y(n26767) );
  OR2X1 U15836 ( .A(n29367), .B(n34113), .Y(n21723) );
  INVX1 U15837 ( .A(n21723), .Y(n26768) );
  OR2X1 U15838 ( .A(n29366), .B(n34100), .Y(n21710) );
  INVX1 U15839 ( .A(n21710), .Y(n26769) );
  OR2X1 U15840 ( .A(n29370), .B(n34152), .Y(n21762) );
  INVX1 U15841 ( .A(n21762), .Y(n26770) );
  INVX1 U15842 ( .A(n21749), .Y(n26771) );
  OR2X1 U15843 ( .A(n29371), .B(n34087), .Y(n21696) );
  INVX1 U15844 ( .A(n21696), .Y(n26772) );
  OR2X1 U15845 ( .A(n29371), .B(n34074), .Y(n21683) );
  INVX1 U15846 ( .A(n21683), .Y(n26773) );
  OR2X1 U15847 ( .A(n29370), .B(n34061), .Y(n21670) );
  INVX1 U15848 ( .A(n21670), .Y(n26774) );
  OR2X1 U15849 ( .A(n29365), .B(n34048), .Y(n21656) );
  INVX1 U15850 ( .A(n21656), .Y(n26775) );
  OR2X1 U15851 ( .A(n29370), .B(n34035), .Y(n21643) );
  INVX1 U15852 ( .A(n21643), .Y(n26776) );
  OR2X1 U15853 ( .A(n29370), .B(n34022), .Y(n21630) );
  INVX1 U15854 ( .A(n21630), .Y(n26777) );
  OR2X1 U15855 ( .A(n29364), .B(n34011), .Y(n21619) );
  INVX1 U15856 ( .A(n21619), .Y(n26778) );
  OR2X1 U15857 ( .A(n29363), .B(n34003), .Y(n21611) );
  INVX1 U15858 ( .A(n21611), .Y(n26779) );
  AND2X2 U15859 ( .A(n30038), .B(n29748), .Y(n29744) );
  AND2X2 U15860 ( .A(n21535), .B(n26781), .Y(n21820) );
  INVX1 U15861 ( .A(n21820), .Y(n26780) );
  AND2X2 U15862 ( .A(n11658), .B(net96578), .Y(n33980) );
  INVX1 U15863 ( .A(n33980), .Y(n26781) );
  INVX8 U15864 ( .A(net96584), .Y(net96578) );
  OR2X1 U15865 ( .A(oc[25]), .B(oc[27]), .Y(n29613) );
  INVX1 U15866 ( .A(n29613), .Y(n26782) );
  BUFX2 U15867 ( .A(n14599), .Y(n26783) );
  BUFX2 U15868 ( .A(n14758), .Y(n26784) );
  BUFX2 U15869 ( .A(n14784), .Y(n26785) );
  BUFX2 U15870 ( .A(n14930), .Y(n26786) );
  BUFX2 U15871 ( .A(n15113), .Y(n26787) );
  AND2X2 U15872 ( .A(n29845), .B(n29728), .Y(n29735) );
  INVX1 U15873 ( .A(n29735), .Y(n26788) );
  AND2X1 U15874 ( .A(n27312), .B(n30457), .Y(n31537) );
  INVX1 U15875 ( .A(n31537), .Y(n26789) );
  AND2X1 U15876 ( .A(n30319), .B(n30440), .Y(n31340) );
  INVX1 U15877 ( .A(n31340), .Y(n26790) );
  AND2X1 U15878 ( .A(n30225), .B(n30418), .Y(n30975) );
  INVX1 U15879 ( .A(n30975), .Y(n26791) );
  AND2X1 U15880 ( .A(n30179), .B(n27323), .Y(n30954) );
  INVX1 U15881 ( .A(n30954), .Y(n26792) );
  AND2X1 U15882 ( .A(n30135), .B(n30426), .Y(n30670) );
  INVX1 U15883 ( .A(n30670), .Y(n26793) );
  AND2X2 U15884 ( .A(n29352), .B(n30562), .Y(n29907) );
  INVX1 U15885 ( .A(n29907), .Y(n26794) );
  AND2X2 U15886 ( .A(n29352), .B(n30601), .Y(n29996) );
  INVX1 U15887 ( .A(n29996), .Y(n26795) );
  AND2X1 U15888 ( .A(n27273), .B(n29821), .Y(n30524) );
  INVX1 U15889 ( .A(n30524), .Y(n26796) );
  AND2X2 U15890 ( .A(n29811), .B(n27314), .Y(n29912) );
  INVX1 U15891 ( .A(n29912), .Y(n26797) );
  INVX1 U15892 ( .A(n29912), .Y(n26798) );
  AND2X2 U15893 ( .A(n29815), .B(n27315), .Y(n30040) );
  INVX1 U15894 ( .A(n30040), .Y(n26799) );
  AND2X1 U15895 ( .A(n27274), .B(n26919), .Y(n16173) );
  INVX1 U15896 ( .A(n16173), .Y(n26800) );
  BUFX2 U15897 ( .A(n16171), .Y(n26801) );
  BUFX2 U15898 ( .A(n16172), .Y(n26802) );
  OR2X1 U15899 ( .A(n34558), .B(n27097), .Y(n16179) );
  AND2X1 U15900 ( .A(n27193), .B(n27101), .Y(n29638) );
  INVX1 U15901 ( .A(n29638), .Y(n26803) );
  AND2X1 U15902 ( .A(n26866), .B(n27187), .Y(n16160) );
  INVX1 U15903 ( .A(n16160), .Y(n26804) );
  AND2X2 U15904 ( .A(n21186), .B(T[3]), .Y(n29656) );
  INVX1 U15905 ( .A(n29656), .Y(n26805) );
  INVX1 U15906 ( .A(n31646), .Y(n26806) );
  INVX1 U15907 ( .A(n31393), .Y(n26807) );
  INVX1 U15908 ( .A(n31024), .Y(n26808) );
  AND2X1 U15909 ( .A(n29221), .B(n27073), .Y(n30785) );
  INVX1 U15910 ( .A(n30785), .Y(n26809) );
  AND2X2 U15911 ( .A(n23301), .B(n29330), .Y(n32792) );
  INVX1 U15912 ( .A(n32792), .Y(n26810) );
  INVX1 U15913 ( .A(n32792), .Y(n26811) );
  INVX1 U15914 ( .A(n29642), .Y(n26812) );
  AND2X2 U15915 ( .A(n30273), .B(n27237), .Y(n32023) );
  INVX1 U15916 ( .A(n32023), .Y(n26813) );
  INVX1 U15917 ( .A(n32023), .Y(n26814) );
  AND2X2 U15918 ( .A(n27265), .B(n30442), .Y(n31933) );
  INVX1 U15919 ( .A(n31933), .Y(n26815) );
  INVX1 U15920 ( .A(n31933), .Y(n26816) );
  AND2X2 U15921 ( .A(n27236), .B(n30458), .Y(n31983) );
  INVX1 U15922 ( .A(n31983), .Y(n26817) );
  INVX1 U15923 ( .A(n31983), .Y(n26818) );
  AND2X2 U15924 ( .A(n29835), .B(n23284), .Y(n33883) );
  INVX1 U15925 ( .A(n33883), .Y(n26819) );
  INVX1 U15926 ( .A(n33883), .Y(n26820) );
  AND2X2 U15927 ( .A(n27322), .B(n29745), .Y(n30012) );
  INVX1 U15928 ( .A(n30012), .Y(n26821) );
  BUFX2 U15929 ( .A(n30023), .Y(n26822) );
  INVX1 U15930 ( .A(n26822), .Y(n29831) );
  OR2X1 U15931 ( .A(n29371), .B(n34164), .Y(n21775) );
  INVX1 U15932 ( .A(n21775), .Y(n26823) );
  OR2X1 U15933 ( .A(n29368), .B(n34125), .Y(n21735) );
  INVX1 U15934 ( .A(n21735), .Y(n26824) );
  OR2X1 U15935 ( .A(n29367), .B(n34112), .Y(n21722) );
  INVX1 U15936 ( .A(n21722), .Y(n26825) );
  OR2X1 U15937 ( .A(n29366), .B(n34099), .Y(n21709) );
  INVX1 U15938 ( .A(n21709), .Y(n26826) );
  OR2X1 U15939 ( .A(n29370), .B(n34151), .Y(n21761) );
  INVX1 U15940 ( .A(n21761), .Y(n26827) );
  INVX1 U15941 ( .A(n21748), .Y(n26828) );
  OR2X1 U15942 ( .A(n29371), .B(n34086), .Y(n21695) );
  INVX1 U15943 ( .A(n21695), .Y(n26829) );
  OR2X1 U15944 ( .A(n29371), .B(n34073), .Y(n21682) );
  INVX1 U15945 ( .A(n21682), .Y(n26830) );
  OR2X1 U15946 ( .A(n29370), .B(n34060), .Y(n21669) );
  INVX1 U15947 ( .A(n21669), .Y(n26831) );
  OR2X1 U15948 ( .A(n29365), .B(n34047), .Y(n21655) );
  INVX1 U15949 ( .A(n21655), .Y(n26832) );
  OR2X1 U15950 ( .A(n29370), .B(n34034), .Y(n21642) );
  INVX1 U15951 ( .A(n21642), .Y(n26833) );
  OR2X1 U15952 ( .A(n29370), .B(n34021), .Y(n21629) );
  INVX1 U15953 ( .A(n21629), .Y(n26834) );
  OR2X1 U15954 ( .A(n29364), .B(n34010), .Y(n21618) );
  INVX1 U15955 ( .A(n21618), .Y(n26835) );
  OR2X1 U15956 ( .A(n29363), .B(n34002), .Y(n21610) );
  INVX1 U15957 ( .A(n21610), .Y(n26836) );
  AND2X2 U15958 ( .A(n29352), .B(n27018), .Y(n30021) );
  INVX1 U15959 ( .A(n30021), .Y(n26837) );
  INVX1 U15960 ( .A(n29605), .Y(n26838) );
  BUFX2 U15961 ( .A(n29548), .Y(n26839) );
  OR2X2 U15962 ( .A(nc[8]), .B(nc[7]), .Y(n29541) );
  INVX1 U15963 ( .A(n29541), .Y(n26840) );
  BUFX2 U15964 ( .A(n14611), .Y(n26841) );
  BUFX2 U15965 ( .A(n14770), .Y(n26842) );
  BUFX2 U15966 ( .A(n14942), .Y(n26843) );
  BUFX2 U15967 ( .A(n14980), .Y(n26844) );
  BUFX2 U15968 ( .A(n15125), .Y(n26845) );
  AND2X1 U15969 ( .A(n27312), .B(n27323), .Y(n31578) );
  INVX1 U15970 ( .A(n31578), .Y(n26846) );
  AND2X1 U15971 ( .A(n30179), .B(n30457), .Y(n30914) );
  INVX1 U15972 ( .A(n30914), .Y(n26847) );
  AND2X2 U15973 ( .A(n29352), .B(n30581), .Y(n29951) );
  INVX1 U15974 ( .A(n29951), .Y(n26848) );
  AND2X2 U15975 ( .A(n29352), .B(n30606), .Y(n30007) );
  INVX1 U15976 ( .A(n30007), .Y(n26849) );
  AND2X1 U15977 ( .A(n27273), .B(n29842), .Y(n30532) );
  INVX1 U15978 ( .A(n30532), .Y(n26850) );
  AND2X1 U15979 ( .A(T[1]), .B(n29689), .Y(n15966) );
  INVX1 U15980 ( .A(n15966), .Y(n26851) );
  AND2X1 U15981 ( .A(n29653), .B(n34351), .Y(n16220) );
  INVX1 U15982 ( .A(n16220), .Y(n26852) );
  AND2X2 U15983 ( .A(n29825), .B(n27314), .Y(n29902) );
  INVX1 U15984 ( .A(n29902), .Y(n26853) );
  BUFX2 U15985 ( .A(n16013), .Y(n26854) );
  AND2X1 U15986 ( .A(n16066), .B(n29674), .Y(n16059) );
  INVX1 U15987 ( .A(n16059), .Y(n26855) );
  AND2X1 U15988 ( .A(T[5]), .B(n16066), .Y(n16060) );
  INVX1 U15989 ( .A(n16060), .Y(n26856) );
  AND2X1 U15990 ( .A(n26928), .B(n27099), .Y(n16007) );
  INVX1 U15991 ( .A(n16007), .Y(n26857) );
  INVX1 U15992 ( .A(n16158), .Y(n26858) );
  BUFX2 U15993 ( .A(n16017), .Y(n26859) );
  AND2X1 U15994 ( .A(n30319), .B(n30418), .Y(n32045) );
  INVX1 U15995 ( .A(n32045), .Y(n26860) );
  AND2X1 U15996 ( .A(n30135), .B(n30432), .Y(n31927) );
  INVX1 U15997 ( .A(n31927), .Y(n26861) );
  INVX1 U15998 ( .A(n31610), .Y(n26862) );
  AND2X1 U15999 ( .A(n29221), .B(n27168), .Y(n31373) );
  INVX1 U16000 ( .A(n31373), .Y(n26863) );
  INVX1 U16001 ( .A(n30987), .Y(n26864) );
  INVX1 U16002 ( .A(n30766), .Y(n26865) );
  AND2X1 U16003 ( .A(T[3]), .B(n26998), .Y(n34591) );
  INVX1 U16004 ( .A(n34591), .Y(n26866) );
  AND2X1 U16005 ( .A(T[4]), .B(n29658), .Y(n16134) );
  INVX1 U16006 ( .A(n16134), .Y(n26867) );
  BUFX2 U16007 ( .A(n15980), .Y(n26868) );
  AND2X2 U16008 ( .A(n23283), .B(n25723), .Y(n32978) );
  INVX1 U16009 ( .A(n32978), .Y(n26869) );
  INVX1 U16010 ( .A(n32978), .Y(n26870) );
  AND2X2 U16011 ( .A(n26271), .B(n34356), .Y(n29643) );
  INVX1 U16012 ( .A(n29643), .Y(n26871) );
  AND2X2 U16013 ( .A(n30227), .B(n27237), .Y(n32000) );
  INVX1 U16014 ( .A(n32000), .Y(n26872) );
  INVX1 U16015 ( .A(n32000), .Y(n26873) );
  AND2X2 U16016 ( .A(n27265), .B(n30476), .Y(n31953) );
  INVX1 U16017 ( .A(n31953), .Y(n26874) );
  INVX1 U16018 ( .A(n31953), .Y(n26875) );
  AND2X2 U16019 ( .A(n27236), .B(n30442), .Y(n31974) );
  INVX1 U16020 ( .A(n31974), .Y(n26876) );
  INVX1 U16021 ( .A(n31974), .Y(n26877) );
  AND2X2 U16022 ( .A(n30626), .B(n30033), .Y(n34218) );
  INVX1 U16023 ( .A(n34218), .Y(n26879) );
  BUFX2 U16024 ( .A(n29989), .Y(n26880) );
  INVX1 U16025 ( .A(n26880), .Y(n29825) );
  OR2X1 U16026 ( .A(n29371), .B(n34163), .Y(n21774) );
  INVX1 U16027 ( .A(n21774), .Y(n26881) );
  OR2X1 U16028 ( .A(n29368), .B(n34124), .Y(n21734) );
  INVX1 U16029 ( .A(n21734), .Y(n26882) );
  OR2X1 U16030 ( .A(n29367), .B(n34111), .Y(n21721) );
  INVX1 U16031 ( .A(n21721), .Y(n26883) );
  OR2X1 U16032 ( .A(n29366), .B(n34098), .Y(n21708) );
  INVX1 U16033 ( .A(n21708), .Y(n26884) );
  OR2X1 U16034 ( .A(n29370), .B(n34150), .Y(n21760) );
  INVX1 U16035 ( .A(n21760), .Y(n26885) );
  INVX1 U16036 ( .A(n21747), .Y(n26886) );
  OR2X1 U16037 ( .A(n29371), .B(n34085), .Y(n21694) );
  INVX1 U16038 ( .A(n21694), .Y(n26887) );
  OR2X1 U16039 ( .A(n29371), .B(n34072), .Y(n21681) );
  INVX1 U16040 ( .A(n21681), .Y(n26888) );
  OR2X1 U16041 ( .A(n29370), .B(n34059), .Y(n21668) );
  INVX1 U16042 ( .A(n21668), .Y(n26889) );
  OR2X1 U16043 ( .A(n29365), .B(n34046), .Y(n21654) );
  INVX1 U16044 ( .A(n21654), .Y(n26890) );
  OR2X1 U16045 ( .A(n29370), .B(n34033), .Y(n21641) );
  INVX1 U16046 ( .A(n21641), .Y(n26891) );
  OR2X1 U16047 ( .A(n29370), .B(n34020), .Y(n21628) );
  INVX1 U16048 ( .A(n21628), .Y(n26892) );
  OR2X1 U16049 ( .A(n29364), .B(n34009), .Y(n21617) );
  INVX1 U16050 ( .A(n21617), .Y(n26893) );
  OR2X1 U16051 ( .A(n29363), .B(n34001), .Y(n21609) );
  INVX1 U16052 ( .A(n21609), .Y(n26894) );
  AND2X2 U16053 ( .A(n31868), .B(n30078), .Y(n31892) );
  AND2X1 U16054 ( .A(net96340), .B(n30629), .Y(n15190) );
  INVX1 U16055 ( .A(n15190), .Y(n26895) );
  INVX1 U16056 ( .A(n29607), .Y(n26896) );
  OR2X1 U16057 ( .A(oc[21]), .B(oc[19]), .Y(n29615) );
  INVX1 U16058 ( .A(n29615), .Y(n26897) );
  AND2X2 U16059 ( .A(n29387), .B(n27103), .Y(n33862) );
  INVX1 U16060 ( .A(n33862), .Y(n26898) );
  AND2X1 U16061 ( .A(n29388), .B(n27191), .Y(n33793) );
  INVX1 U16062 ( .A(n33793), .Y(n26899) );
  AND2X2 U16063 ( .A(n29416), .B(n21375), .Y(n33833) );
  INVX1 U16064 ( .A(n33833), .Y(n26900) );
  OR2X2 U16065 ( .A(nc[23]), .B(nc[22]), .Y(n29529) );
  INVX1 U16066 ( .A(n29529), .Y(n26901) );
  BUFX2 U16067 ( .A(n14623), .Y(n26902) );
  BUFX2 U16068 ( .A(n14808), .Y(n26903) );
  BUFX2 U16069 ( .A(n14882), .Y(n26904) );
  BUFX2 U16070 ( .A(n14992), .Y(n26905) );
  BUFX2 U16071 ( .A(n15137), .Y(n26906) );
  AND2X2 U16072 ( .A(n29352), .B(n30494), .Y(n29765) );
  INVX1 U16073 ( .A(n29765), .Y(n26907) );
  AND2X1 U16074 ( .A(n30426), .B(n27324), .Y(n31776) );
  INVX1 U16075 ( .A(n31776), .Y(n26908) );
  AND2X1 U16076 ( .A(n30409), .B(n30440), .Y(n31660) );
  INVX1 U16077 ( .A(n31660), .Y(n26909) );
  AND2X1 U16078 ( .A(n30272), .B(n30457), .Y(n31233) );
  INVX1 U16079 ( .A(n31233), .Y(n26910) );
  AND2X1 U16080 ( .A(n30225), .B(n27323), .Y(n31116) );
  INVX1 U16081 ( .A(n31116), .Y(n26911) );
  AND2X2 U16082 ( .A(n29352), .B(n30566), .Y(n29917) );
  INVX1 U16083 ( .A(n29917), .Y(n26912) );
  AND2X1 U16084 ( .A(n27273), .B(n29860), .Y(n30542) );
  INVX1 U16085 ( .A(n30542), .Y(n26913) );
  AND2X1 U16086 ( .A(n29681), .B(n34351), .Y(n15988) );
  INVX1 U16087 ( .A(n15988), .Y(n26914) );
  BUFX2 U16088 ( .A(n16014), .Y(n26915) );
  OR2X1 U16089 ( .A(n34564), .B(n27006), .Y(n16021) );
  AND2X2 U16090 ( .A(n27314), .B(n29967), .Y(n29968) );
  INVX1 U16091 ( .A(n29968), .Y(n26916) );
  INVX1 U16092 ( .A(n15932), .Y(n26917) );
  AND2X1 U16093 ( .A(n27197), .B(n27100), .Y(n16157) );
  INVX1 U16094 ( .A(n16157), .Y(n26918) );
  BUFX2 U16095 ( .A(n16175), .Y(n26919) );
  BUFX2 U16096 ( .A(n16204), .Y(n26920) );
  AND2X1 U16097 ( .A(n30179), .B(n30449), .Y(n31977) );
  INVX1 U16098 ( .A(n31977), .Y(n26921) );
  INVX1 U16099 ( .A(n31591), .Y(n26922) );
  INVX1 U16100 ( .A(n31353), .Y(n26923) );
  AND2X1 U16101 ( .A(n29221), .B(n26992), .Y(n30946) );
  INVX1 U16102 ( .A(n30946), .Y(n26924) );
  AND2X1 U16103 ( .A(n29221), .B(n26993), .Y(n30745) );
  INVX1 U16104 ( .A(n30745), .Y(n26925) );
  AND2X1 U16105 ( .A(n27312), .B(n30432), .Y(n32084) );
  INVX1 U16106 ( .A(n32084), .Y(n26926) );
  AND2X1 U16107 ( .A(n30319), .B(n27311), .Y(n32068) );
  INVX1 U16108 ( .A(n32068), .Y(n26927) );
  AND2X1 U16109 ( .A(n29673), .B(T[3]), .Y(n34594) );
  INVX1 U16110 ( .A(n34594), .Y(n26928) );
  AND2X1 U16111 ( .A(T[4]), .B(n29650), .Y(n16215) );
  INVX1 U16112 ( .A(n16215), .Y(n26929) );
  AND2X1 U16113 ( .A(n29688), .B(n34372), .Y(n15964) );
  INVX1 U16114 ( .A(n15964), .Y(n26930) );
  AND2X2 U16115 ( .A(n23298), .B(n29331), .Y(n32988) );
  INVX1 U16116 ( .A(n32988), .Y(n26931) );
  AND2X2 U16117 ( .A(n29748), .B(n27018), .Y(n29891) );
  INVX1 U16118 ( .A(n29891), .Y(n26932) );
  AND2X1 U16119 ( .A(n29659), .B(n34356), .Y(n16132) );
  INVX1 U16120 ( .A(n16132), .Y(n26933) );
  AND2X2 U16121 ( .A(n27265), .B(n27237), .Y(n31923) );
  INVX1 U16122 ( .A(n31923), .Y(n26934) );
  INVX1 U16123 ( .A(n31923), .Y(n26935) );
  AND2X2 U16124 ( .A(n27236), .B(n30433), .Y(n31969) );
  INVX1 U16125 ( .A(n31969), .Y(n26936) );
  INVX1 U16126 ( .A(n31969), .Y(n26937) );
  AND2X2 U16127 ( .A(n21183), .B(n34360), .Y(n29655) );
  INVX1 U16128 ( .A(n29655), .Y(n26938) );
  BUFX2 U16129 ( .A(n29956), .Y(n26939) );
  INVX1 U16130 ( .A(n33617), .Y(n26940) );
  AND2X2 U16131 ( .A(n29835), .B(n27303), .Y(n33704) );
  INVX1 U16132 ( .A(n33704), .Y(n26941) );
  INVX1 U16133 ( .A(n33704), .Y(n26942) );
  AND2X2 U16134 ( .A(n30442), .B(n30475), .Y(n32141) );
  INVX4 U16135 ( .A(n32141), .Y(n26943) );
  AND2X2 U16136 ( .A(n30411), .B(n30458), .Y(n32124) );
  INVX4 U16137 ( .A(n32124), .Y(n26944) );
  AND2X2 U16138 ( .A(n30273), .B(n30476), .Y(n32041) );
  INVX1 U16139 ( .A(n32041), .Y(n26945) );
  INVX1 U16140 ( .A(n32041), .Y(n26946) );
  INVX1 U16141 ( .A(n32041), .Y(n26947) );
  AND2X2 U16142 ( .A(n27248), .B(n27315), .Y(n30035) );
  INVX1 U16143 ( .A(n30035), .Y(n26948) );
  INVX2 U16144 ( .A(n33933), .Y(n33934) );
  OR2X1 U16145 ( .A(n29371), .B(n34162), .Y(n21773) );
  INVX1 U16146 ( .A(n21773), .Y(n26950) );
  OR2X1 U16147 ( .A(n29368), .B(n34123), .Y(n21733) );
  INVX1 U16148 ( .A(n21733), .Y(n26951) );
  OR2X1 U16149 ( .A(n29367), .B(n34110), .Y(n21720) );
  INVX1 U16150 ( .A(n21720), .Y(n26952) );
  OR2X1 U16151 ( .A(n29366), .B(n34097), .Y(n21707) );
  INVX1 U16152 ( .A(n21707), .Y(n26953) );
  OR2X1 U16153 ( .A(n29370), .B(n34149), .Y(n21759) );
  INVX1 U16154 ( .A(n21759), .Y(n26954) );
  INVX1 U16155 ( .A(n21746), .Y(n26955) );
  OR2X1 U16156 ( .A(n29371), .B(n34084), .Y(n21693) );
  INVX1 U16157 ( .A(n21693), .Y(n26956) );
  OR2X1 U16158 ( .A(n29371), .B(n34071), .Y(n21680) );
  INVX1 U16159 ( .A(n21680), .Y(n26957) );
  OR2X1 U16160 ( .A(n29370), .B(n34058), .Y(n21667) );
  INVX1 U16161 ( .A(n21667), .Y(n26958) );
  OR2X1 U16162 ( .A(n29365), .B(n34045), .Y(n21653) );
  INVX1 U16163 ( .A(n21653), .Y(n26959) );
  OR2X1 U16164 ( .A(n29371), .B(n34032), .Y(n21640) );
  INVX1 U16165 ( .A(n21640), .Y(n26960) );
  OR2X1 U16166 ( .A(n29370), .B(n34019), .Y(n21627) );
  INVX1 U16167 ( .A(n21627), .Y(n26961) );
  OR2X1 U16168 ( .A(n29364), .B(n34005), .Y(n21613) );
  INVX1 U16169 ( .A(n21613), .Y(n26962) );
  OR2X1 U16170 ( .A(n29363), .B(n34000), .Y(n21608) );
  INVX1 U16171 ( .A(n21608), .Y(n26963) );
  AND2X2 U16172 ( .A(n29381), .B(n30474), .Y(n30631) );
  AND2X2 U16173 ( .A(n29389), .B(n27207), .Y(n33662) );
  INVX1 U16174 ( .A(n33662), .Y(n26964) );
  INVX4 U16175 ( .A(n29392), .Y(n29389) );
  AND2X2 U16176 ( .A(n29416), .B(n27103), .Y(n33856) );
  INVX1 U16177 ( .A(n33856), .Y(n26965) );
  BUFX2 U16178 ( .A(n14647), .Y(n26966) );
  BUFX2 U16179 ( .A(n14686), .Y(n26967) );
  BUFX2 U16180 ( .A(n14820), .Y(n26968) );
  BUFX2 U16181 ( .A(n14966), .Y(n26969) );
  BUFX2 U16182 ( .A(n15149), .Y(n26970) );
  INVX2 U16183 ( .A(n3773), .Y(n34230) );
  AND2X1 U16184 ( .A(n31770), .B(net96340), .Y(n31777) );
  INVX1 U16185 ( .A(n31777), .Y(n26971) );
  AND2X1 U16186 ( .A(n31070), .B(net96340), .Y(n31077) );
  INVX1 U16187 ( .A(n31077), .Y(n26972) );
  AND2X1 U16188 ( .A(n31187), .B(net96340), .Y(n31194) );
  INVX1 U16189 ( .A(n31194), .Y(n26973) );
  AND2X1 U16190 ( .A(n30440), .B(n27324), .Y(n31815) );
  INVX1 U16191 ( .A(n31815), .Y(n26974) );
  AND2X1 U16192 ( .A(n30409), .B(n30426), .Y(n31624) );
  INVX1 U16193 ( .A(n31624), .Y(n26975) );
  AND2X1 U16194 ( .A(n30272), .B(n27323), .Y(n31273) );
  INVX1 U16195 ( .A(n31273), .Y(n26976) );
  AND2X1 U16196 ( .A(n30225), .B(n30457), .Y(n31076) );
  INVX1 U16197 ( .A(n31076), .Y(n26977) );
  AND2X2 U16198 ( .A(n29352), .B(n30591), .Y(n29973) );
  INVX1 U16199 ( .A(n29973), .Y(n26979) );
  INVX1 U16200 ( .A(n30496), .Y(n26980) );
  INVX1 U16201 ( .A(n29767), .Y(n26981) );
  AND2X2 U16202 ( .A(n27115), .B(n27204), .Y(n29766) );
  INVX1 U16203 ( .A(n29766), .Y(n26982) );
  INVX1 U16204 ( .A(net108311), .Y(net104600) );
  AND2X2 U16205 ( .A(n29815), .B(n27314), .Y(n29943) );
  INVX1 U16206 ( .A(n29943), .Y(n26983) );
  AND2X2 U16207 ( .A(n29811), .B(n27315), .Y(n30002) );
  INVX1 U16208 ( .A(n30002), .Y(n26984) );
  INVX1 U16209 ( .A(n14478), .Y(n26985) );
  OR2X2 U16210 ( .A(n21137), .B(n23204), .Y(n29620) );
  INVX1 U16211 ( .A(n29620), .Y(n26986) );
  AND2X1 U16212 ( .A(n29221), .B(n27167), .Y(n31570) );
  INVX1 U16213 ( .A(n31570), .Y(n26987) );
  AND2X1 U16214 ( .A(n29221), .B(n27071), .Y(n31333) );
  INVX1 U16215 ( .A(n31333), .Y(n26988) );
  INVX1 U16216 ( .A(n30967), .Y(n26989) );
  INVX1 U16217 ( .A(n30726), .Y(n26990) );
  AND2X1 U16218 ( .A(n27312), .B(n30418), .Y(n32076) );
  INVX1 U16219 ( .A(n32076), .Y(n26991) );
  AND2X1 U16220 ( .A(n30179), .B(n27311), .Y(n31987) );
  INVX1 U16221 ( .A(n31987), .Y(n26992) );
  AND2X1 U16222 ( .A(n30135), .B(n30449), .Y(n31937) );
  INVX1 U16223 ( .A(n31937), .Y(n26993) );
  AND2X1 U16224 ( .A(n29686), .B(n34385), .Y(n15971) );
  INVX1 U16225 ( .A(n15971), .Y(n26994) );
  AND2X1 U16226 ( .A(T[4]), .B(n29675), .Y(n15983) );
  INVX1 U16227 ( .A(n15983), .Y(n26995) );
  AND2X2 U16228 ( .A(n23299), .B(n29330), .Y(n32882) );
  INVX1 U16229 ( .A(n21188), .Y(n26996) );
  AND2X2 U16230 ( .A(n27191), .B(n27121), .Y(n30504) );
  INVX1 U16231 ( .A(n30504), .Y(n26997) );
  AND2X2 U16232 ( .A(n20977), .B(n25722), .Y(n29652) );
  INVX1 U16233 ( .A(n29652), .Y(n26998) );
  AND2X1 U16234 ( .A(T[0]), .B(n27098), .Y(n34572) );
  INVX1 U16235 ( .A(n34572), .Y(n26999) );
  AND2X1 U16236 ( .A(n29671), .B(n34356), .Y(n16055) );
  INVX1 U16237 ( .A(n16055), .Y(n27000) );
  AND2X2 U16238 ( .A(n27265), .B(n30464), .Y(n31948) );
  INVX1 U16239 ( .A(n31948), .Y(n27001) );
  INVX1 U16240 ( .A(n31948), .Y(n27002) );
  AND2X2 U16241 ( .A(n27236), .B(n30450), .Y(n31978) );
  INVX1 U16242 ( .A(n31978), .Y(n27003) );
  INVX1 U16243 ( .A(n31978), .Y(n27004) );
  INVX1 U16244 ( .A(n16184), .Y(n27005) );
  BUFX2 U16245 ( .A(n16012), .Y(n27006) );
  BUFX2 U16246 ( .A(n16167), .Y(n27007) );
  AND2X1 U16247 ( .A(n29680), .B(n34360), .Y(n15953) );
  INVX1 U16248 ( .A(n15953), .Y(n27008) );
  AND2X2 U16249 ( .A(n30411), .B(n30442), .Y(n32118) );
  INVX4 U16250 ( .A(n32118), .Y(n27009) );
  AND2X2 U16251 ( .A(n30273), .B(n30458), .Y(n32035) );
  INVX1 U16252 ( .A(n32035), .Y(n27010) );
  INVX1 U16253 ( .A(n32035), .Y(n27011) );
  INVX1 U16254 ( .A(n32035), .Y(n27012) );
  AND2X2 U16255 ( .A(n30227), .B(n30476), .Y(n32017) );
  INVX1 U16256 ( .A(n32017), .Y(n27013) );
  INVX1 U16257 ( .A(n32017), .Y(n27014) );
  INVX1 U16258 ( .A(n32017), .Y(n27015) );
  BUFX2 U16259 ( .A(n30001), .Y(n27016) );
  INVX1 U16260 ( .A(n27016), .Y(n29811) );
  BUFX2 U16261 ( .A(n30036), .Y(n27017) );
  INVX1 U16262 ( .A(n27017), .Y(n29815) );
  AND2X2 U16263 ( .A(n25170), .B(n29633), .Y(n30073) );
  INVX1 U16264 ( .A(n21055), .Y(n27018) );
  AND2X2 U16265 ( .A(n29835), .B(n25749), .Y(n33814) );
  INVX1 U16266 ( .A(n33814), .Y(n27020) );
  INVX1 U16267 ( .A(n33814), .Y(n27021) );
  INVX1 U16268 ( .A(n27020), .Y(n33829) );
  AND2X2 U16269 ( .A(n29968), .B(n21106), .Y(n32855) );
  INVX1 U16270 ( .A(n32855), .Y(n27022) );
  INVX1 U16271 ( .A(n32855), .Y(n27023) );
  INVX1 U16272 ( .A(n32855), .Y(n27024) );
  BUFX2 U16273 ( .A(net95456), .Y(net104480) );
  AND2X2 U16274 ( .A(n30033), .B(n21106), .Y(n32945) );
  INVX1 U16275 ( .A(n32945), .Y(n27025) );
  INVX1 U16276 ( .A(n32945), .Y(n27026) );
  INVX1 U16277 ( .A(n32945), .Y(n27027) );
  OR2X1 U16278 ( .A(n29371), .B(n34161), .Y(n21772) );
  INVX1 U16279 ( .A(n21772), .Y(n27028) );
  OR2X1 U16280 ( .A(n29368), .B(n34122), .Y(n21732) );
  INVX1 U16281 ( .A(n21732), .Y(n27029) );
  OR2X1 U16282 ( .A(n29367), .B(n34109), .Y(n21719) );
  INVX1 U16283 ( .A(n21719), .Y(n27030) );
  OR2X1 U16284 ( .A(n29366), .B(n34096), .Y(n21706) );
  INVX1 U16285 ( .A(n21706), .Y(n27031) );
  OR2X1 U16286 ( .A(n29370), .B(n34148), .Y(n21758) );
  INVX1 U16287 ( .A(n21758), .Y(n27032) );
  INVX1 U16288 ( .A(n21745), .Y(n27033) );
  OR2X1 U16289 ( .A(n29371), .B(n34083), .Y(n21692) );
  INVX1 U16290 ( .A(n21692), .Y(n27034) );
  OR2X1 U16291 ( .A(n29370), .B(n34070), .Y(n21679) );
  INVX1 U16292 ( .A(n21679), .Y(n27035) );
  OR2X1 U16293 ( .A(n29370), .B(n34057), .Y(n21665) );
  INVX1 U16294 ( .A(n21665), .Y(n27036) );
  OR2X1 U16295 ( .A(n29365), .B(n34044), .Y(n21652) );
  INVX1 U16296 ( .A(n21652), .Y(n27037) );
  OR2X1 U16297 ( .A(n29370), .B(n34031), .Y(n21639) );
  INVX1 U16298 ( .A(n21639), .Y(n27038) );
  OR2X1 U16299 ( .A(n29370), .B(n34018), .Y(n21626) );
  INVX1 U16300 ( .A(n21626), .Y(n27039) );
  OR2X1 U16301 ( .A(n29364), .B(n34004), .Y(n21612) );
  INVX1 U16302 ( .A(n21612), .Y(n27040) );
  OR2X1 U16303 ( .A(n29363), .B(n33997), .Y(n21605) );
  INVX1 U16304 ( .A(n21605), .Y(n27041) );
  AND2X2 U16305 ( .A(n29416), .B(n27191), .Y(n33788) );
  INVX1 U16306 ( .A(n33788), .Y(n27045) );
  INVX4 U16307 ( .A(n29418), .Y(n29416) );
  AND2X2 U16308 ( .A(n29415), .B(n21378), .Y(n33766) );
  INVX1 U16309 ( .A(n33766), .Y(n27046) );
  AND2X2 U16310 ( .A(n29415), .B(n27207), .Y(n33657) );
  INVX1 U16311 ( .A(n33657), .Y(n27047) );
  INVX4 U16312 ( .A(n29418), .Y(n29415) );
  OR2X2 U16313 ( .A(n32587), .B(n21155), .Y(n32588) );
  INVX1 U16314 ( .A(n32588), .Y(n27048) );
  BUFX2 U16315 ( .A(n30650), .Y(n29207) );
  BUFX2 U16316 ( .A(n14587), .Y(n27049) );
  BUFX2 U16317 ( .A(n14698), .Y(n27050) );
  BUFX2 U16318 ( .A(n14844), .Y(n27051) );
  BUFX2 U16319 ( .A(n14954), .Y(n27052) );
  BUFX2 U16320 ( .A(n15064), .Y(n27053) );
  AND2X1 U16321 ( .A(n30457), .B(n27324), .Y(n31855) );
  INVX1 U16322 ( .A(n31855), .Y(n27054) );
  AND2X1 U16323 ( .A(n30409), .B(n27323), .Y(n31738) );
  INVX1 U16324 ( .A(n31738), .Y(n27055) );
  AND2X1 U16325 ( .A(n30272), .B(n30426), .Y(n31156) );
  INVX1 U16326 ( .A(n31156), .Y(n27056) );
  AND2X1 U16327 ( .A(n30225), .B(n30440), .Y(n31038) );
  INVX1 U16328 ( .A(n31038), .Y(n27057) );
  INVX1 U16329 ( .A(n23206), .Y(n27058) );
  AND2X2 U16330 ( .A(n29713), .B(n29946), .Y(n29726) );
  INVX1 U16331 ( .A(n29726), .Y(n27059) );
  BUFX2 U16332 ( .A(n15940), .Y(n27060) );
  OR2X1 U16333 ( .A(n34569), .B(n27185), .Y(n15947) );
  AND2X2 U16334 ( .A(n27294), .B(n29967), .Y(n29807) );
  INVX1 U16335 ( .A(n29807), .Y(n27061) );
  AND2X2 U16336 ( .A(net137830), .B(Setup[1]), .Y(n30482) );
  INVX1 U16337 ( .A(n30482), .Y(n27062) );
  OR2X2 U16338 ( .A(address[3]), .B(n27192), .Y(n14576) );
  INVX1 U16339 ( .A(n14576), .Y(n27063) );
  AND2X2 U16340 ( .A(net95156), .B(net108803), .Y(n29698) );
  INVX1 U16341 ( .A(n29698), .Y(n27064) );
  INVX1 U16342 ( .A(n29698), .Y(n27065) );
  AND2X1 U16343 ( .A(n27312), .B(n30449), .Y(n32091) );
  INVX1 U16344 ( .A(n32091), .Y(n27066) );
  INVX1 U16345 ( .A(n31550), .Y(n27067) );
  INVX1 U16346 ( .A(n31315), .Y(n27068) );
  INVX1 U16347 ( .A(n30927), .Y(n27069) );
  INVX1 U16348 ( .A(n30706), .Y(n27070) );
  AND2X1 U16349 ( .A(n30319), .B(n30432), .Y(n32053) );
  INVX1 U16350 ( .A(n32053), .Y(n27071) );
  AND2X1 U16351 ( .A(n30179), .B(n30418), .Y(n31958) );
  INVX1 U16352 ( .A(n31958), .Y(n27072) );
  AND2X1 U16353 ( .A(n30135), .B(n27311), .Y(n31947) );
  INVX1 U16354 ( .A(n31947), .Y(n27073) );
  INVX1 U16355 ( .A(n34320), .Y(n27074) );
  AND2X2 U16356 ( .A(n30186), .B(n29672), .Y(n29674) );
  INVX1 U16357 ( .A(n29674), .Y(n27075) );
  AND2X1 U16358 ( .A(T[4]), .B(n29669), .Y(n16057) );
  INVX1 U16359 ( .A(n16057), .Y(n27076) );
  AND2X1 U16360 ( .A(n29666), .B(n34372), .Y(n16115) );
  INVX1 U16361 ( .A(n16115), .Y(n27077) );
  AND2X2 U16362 ( .A(n23286), .B(n29330), .Y(n32871) );
  INVX1 U16363 ( .A(n32871), .Y(n27078) );
  AND2X2 U16364 ( .A(n21375), .B(n27206), .Y(n30495) );
  INVX1 U16365 ( .A(n30495), .Y(n27079) );
  AND2X2 U16366 ( .A(n23296), .B(n21106), .Y(n29794) );
  INVX1 U16367 ( .A(n29794), .Y(n27080) );
  AND2X2 U16368 ( .A(n21224), .B(n27322), .Y(n29967) );
  INVX1 U16369 ( .A(n29967), .Y(n27081) );
  INVX1 U16370 ( .A(n29967), .Y(n27082) );
  AND2X2 U16371 ( .A(n27302), .B(n29465), .Y(n29477) );
  INVX1 U16372 ( .A(n29477), .Y(n27083) );
  AND2X2 U16373 ( .A(n26073), .B(alt5_net95676), .Y(n27302) );
  AND2X1 U16374 ( .A(n29648), .B(n29647), .Y(n34597) );
  INVX1 U16375 ( .A(n34597), .Y(n27085) );
  AND2X1 U16376 ( .A(n29651), .B(n34356), .Y(n16213) );
  INVX1 U16377 ( .A(n16213), .Y(n27086) );
  AND2X2 U16378 ( .A(n27265), .B(n30450), .Y(n31938) );
  INVX1 U16379 ( .A(n31938), .Y(n27087) );
  INVX1 U16380 ( .A(n31938), .Y(n27088) );
  AND2X2 U16381 ( .A(n27265), .B(n30433), .Y(n31928) );
  INVX1 U16382 ( .A(n31928), .Y(n27089) );
  INVX1 U16383 ( .A(n31928), .Y(n27090) );
  AND2X2 U16384 ( .A(n27245), .B(n29461), .Y(n27265) );
  AND2X2 U16385 ( .A(n27236), .B(n30476), .Y(n31994) );
  INVX1 U16386 ( .A(n31994), .Y(n27091) );
  INVX1 U16387 ( .A(n31994), .Y(n27092) );
  AND2X2 U16388 ( .A(n27236), .B(n30464), .Y(n31988) );
  INVX1 U16389 ( .A(n31988), .Y(n27093) );
  INVX1 U16390 ( .A(n31988), .Y(n27094) );
  AND2X2 U16391 ( .A(n27245), .B(n28606), .Y(n27236) );
  INVX1 U16392 ( .A(n16103), .Y(n27095) );
  INVX1 U16393 ( .A(n15952), .Y(n27096) );
  BUFX2 U16394 ( .A(n16170), .Y(n27097) );
  AND2X2 U16395 ( .A(n30127), .B(n31917), .Y(n29687) );
  INVX1 U16396 ( .A(n29687), .Y(n27098) );
  INVX1 U16397 ( .A(n16027), .Y(n27099) );
  AND2X2 U16398 ( .A(n21007), .B(n34379), .Y(n16187) );
  INVX1 U16399 ( .A(n16187), .Y(n27100) );
  AND2X2 U16400 ( .A(n29683), .B(T[1]), .Y(n16198) );
  INVX1 U16401 ( .A(n16198), .Y(n27101) );
  AND2X2 U16402 ( .A(n29835), .B(n29968), .Y(n33860) );
  INVX1 U16403 ( .A(n33860), .Y(n27102) );
  INVX1 U16404 ( .A(n33860), .Y(n27103) );
  AND2X2 U16405 ( .A(n27237), .B(n30475), .Y(n32135) );
  INVX1 U16406 ( .A(n32135), .Y(n27104) );
  INVX1 U16407 ( .A(n32135), .Y(n27105) );
  INVX1 U16408 ( .A(n32135), .Y(n27106) );
  AND2X2 U16409 ( .A(n27272), .B(n26144), .Y(n27237) );
  AND2X2 U16410 ( .A(n30273), .B(n30442), .Y(n32029) );
  INVX1 U16411 ( .A(n32029), .Y(n27107) );
  INVX1 U16412 ( .A(n32029), .Y(n27108) );
  INVX1 U16413 ( .A(n32029), .Y(n27109) );
  AND2X2 U16414 ( .A(n30227), .B(n30458), .Y(n32011) );
  INVX1 U16415 ( .A(n32011), .Y(n27110) );
  INVX1 U16416 ( .A(n32011), .Y(n27111) );
  INVX1 U16417 ( .A(n32011), .Y(n27112) );
  AND2X2 U16418 ( .A(n23441), .B(n34385), .Y(n16203) );
  INVX1 U16419 ( .A(n16203), .Y(n27113) );
  AND2X2 U16420 ( .A(states[1]), .B(n29527), .Y(n30078) );
  AND2X2 U16421 ( .A(n34498), .B(net109585), .Y(n30038) );
  INVX1 U16422 ( .A(n30038), .Y(n27114) );
  AND2X2 U16423 ( .A(n23288), .B(n29331), .Y(n32991) );
  INVX4 U16424 ( .A(n32991), .Y(n27115) );
  AND2X2 U16425 ( .A(n27248), .B(n27313), .Y(n29879) );
  INVX1 U16426 ( .A(n29879), .Y(n27116) );
  INVX1 U16427 ( .A(n32185), .Y(n27117) );
  INVX1 U16428 ( .A(n32185), .Y(n27118) );
  AND2X2 U16429 ( .A(n23294), .B(n21106), .Y(n32950) );
  INVX1 U16430 ( .A(n32950), .Y(n27119) );
  INVX1 U16431 ( .A(n32950), .Y(n27120) );
  INVX1 U16432 ( .A(n32950), .Y(n27121) );
  OR2X1 U16433 ( .A(reset), .B(Setup[0]), .Y(n21324) );
  INVX2 U16434 ( .A(n21324), .Y(n27122) );
  OR2X1 U16435 ( .A(n29371), .B(n34160), .Y(n21771) );
  INVX1 U16436 ( .A(n21771), .Y(n27123) );
  OR2X1 U16437 ( .A(n29368), .B(n34121), .Y(n21731) );
  INVX1 U16438 ( .A(n21731), .Y(n27124) );
  OR2X1 U16439 ( .A(n29367), .B(n34108), .Y(n21718) );
  INVX1 U16440 ( .A(n21718), .Y(n27125) );
  OR2X1 U16441 ( .A(n29366), .B(n34095), .Y(n21705) );
  INVX1 U16442 ( .A(n21705), .Y(n27126) );
  OR2X1 U16443 ( .A(n29370), .B(n34147), .Y(n21757) );
  INVX1 U16444 ( .A(n21757), .Y(n27127) );
  INVX1 U16445 ( .A(n21744), .Y(n27128) );
  OR2X1 U16446 ( .A(n29371), .B(n34082), .Y(n21691) );
  INVX1 U16447 ( .A(n21691), .Y(n27129) );
  OR2X1 U16448 ( .A(n29370), .B(n34069), .Y(n21678) );
  INVX1 U16449 ( .A(n21678), .Y(n27130) );
  OR2X1 U16450 ( .A(n29370), .B(n34056), .Y(n21664) );
  INVX1 U16451 ( .A(n21664), .Y(n27131) );
  OR2X1 U16452 ( .A(n29365), .B(n34043), .Y(n21651) );
  INVX1 U16453 ( .A(n21651), .Y(n27132) );
  OR2X1 U16454 ( .A(n29370), .B(n34030), .Y(n21638) );
  INVX1 U16455 ( .A(n21638), .Y(n27133) );
  OR2X1 U16456 ( .A(n29370), .B(n34017), .Y(n21625) );
  INVX1 U16457 ( .A(n21625), .Y(n27134) );
  OR2X2 U16458 ( .A(n29364), .B(n34008), .Y(n21616) );
  INVX1 U16459 ( .A(n21616), .Y(n27135) );
  OR2X2 U16460 ( .A(n29364), .B(n34007), .Y(n21615) );
  INVX1 U16461 ( .A(n21615), .Y(n27136) );
  INVX4 U16462 ( .A(n29378), .Y(n29364) );
  OR2X2 U16463 ( .A(n29364), .B(n34006), .Y(n21614) );
  INVX1 U16464 ( .A(n21614), .Y(n27137) );
  OR2X2 U16465 ( .A(n29363), .B(n33999), .Y(n21607) );
  INVX1 U16466 ( .A(n21607), .Y(n27138) );
  OR2X2 U16467 ( .A(n29363), .B(n33998), .Y(n21606) );
  INVX1 U16468 ( .A(n21606), .Y(n27139) );
  INVX4 U16469 ( .A(n29377), .Y(n29363) );
  AND2X2 U16470 ( .A(n29381), .B(n29196), .Y(n30636) );
  AND2X2 U16471 ( .A(n29241), .B(n31868), .Y(n31862) );
  INVX1 U16472 ( .A(n31862), .Y(n27146) );
  AND2X2 U16473 ( .A(net90053), .B(net96340), .Y(n34224) );
  INVX1 U16474 ( .A(n34224), .Y(n27147) );
  BUFX2 U16475 ( .A(n14448), .Y(n27148) );
  BUFX2 U16476 ( .A(n14561), .Y(n27149) );
  BUFX2 U16477 ( .A(n15016), .Y(n27150) );
  BUFX2 U16478 ( .A(n15167), .Y(n27151) );
  AND2X2 U16479 ( .A(n27247), .B(n29321), .Y(n31922) );
  INVX1 U16480 ( .A(n31922), .Y(n27152) );
  AND2X2 U16481 ( .A(Setup[1]), .B(n29703), .Y(n29704) );
  INVX1 U16482 ( .A(n29704), .Y(n27153) );
  AND2X1 U16483 ( .A(n30409), .B(n30457), .Y(n31698) );
  INVX1 U16484 ( .A(n31698), .Y(n27154) );
  AND2X1 U16485 ( .A(n30272), .B(n30440), .Y(n31193) );
  INVX1 U16486 ( .A(n31193), .Y(n27155) );
  AND2X1 U16487 ( .A(n30225), .B(n30426), .Y(n31001) );
  INVX1 U16488 ( .A(n31001), .Y(n27156) );
  AND2X1 U16489 ( .A(n30327), .B(n30126), .Y(n31914) );
  INVX1 U16490 ( .A(n31914), .Y(n27157) );
  AND2X1 U16491 ( .A(n34352), .B(n34351), .Y(n34366) );
  INVX1 U16492 ( .A(n34366), .Y(n27158) );
  BUFX2 U16493 ( .A(n33176), .Y(n27159) );
  INVX2 U16494 ( .A(n3772), .Y(n34280) );
  AND2X2 U16495 ( .A(n29683), .B(n21007), .Y(n30086) );
  INVX1 U16496 ( .A(n30086), .Y(n27160) );
  INVX1 U16497 ( .A(n29561), .Y(n33928) );
  AND2X1 U16498 ( .A(n27273), .B(n29868), .Y(n30547) );
  INVX1 U16499 ( .A(n30547), .Y(n27161) );
  AND2X2 U16500 ( .A(n21217), .B(n26339), .Y(n29679) );
  INVX1 U16501 ( .A(n29679), .Y(n27162) );
  INVX1 U16502 ( .A(n29593), .Y(n34203) );
  INVX1 U16503 ( .A(n31530), .Y(n27163) );
  INVX1 U16504 ( .A(n31296), .Y(n27164) );
  INVX1 U16505 ( .A(n30906), .Y(n27165) );
  INVX1 U16506 ( .A(n30683), .Y(n27166) );
  AND2X1 U16507 ( .A(n27312), .B(n27311), .Y(n32100) );
  INVX1 U16508 ( .A(n32100), .Y(n27167) );
  AND2X1 U16509 ( .A(n30319), .B(n30449), .Y(n32060) );
  INVX1 U16510 ( .A(n32060), .Y(n27168) );
  AND2X1 U16511 ( .A(n30179), .B(n30432), .Y(n31968) );
  INVX1 U16512 ( .A(n31968), .Y(n27169) );
  AND2X1 U16513 ( .A(n30135), .B(n30418), .Y(n31916) );
  INVX1 U16514 ( .A(n31916), .Y(n27170) );
  AND2X2 U16515 ( .A(n30186), .B(n25205), .Y(n29661) );
  INVX1 U16516 ( .A(n29661), .Y(n27171) );
  AND2X2 U16517 ( .A(n25167), .B(n21560), .Y(n33079) );
  BUFX2 U16518 ( .A(n34213), .Y(n27173) );
  AND2X2 U16519 ( .A(n21378), .B(n27080), .Y(n30509) );
  INVX1 U16520 ( .A(n30509), .Y(n27174) );
  AND2X2 U16521 ( .A(n34189), .B(n27257), .Y(n29685) );
  INVX1 U16522 ( .A(n29685), .Y(n27176) );
  AND2X1 U16523 ( .A(n29677), .B(n34356), .Y(n15981) );
  INVX1 U16524 ( .A(n15981), .Y(n27177) );
  AND2X1 U16525 ( .A(n27323), .B(n27324), .Y(n32461) );
  INVX1 U16526 ( .A(n32461), .Y(n27179) );
  AND2X2 U16527 ( .A(n29207), .B(n25334), .Y(n13709) );
  INVX1 U16528 ( .A(n13709), .Y(n27180) );
  INVX1 U16529 ( .A(n13709), .Y(n27181) );
  INVX1 U16530 ( .A(n27180), .Y(n29579) );
  INVX1 U16531 ( .A(n16026), .Y(n27182) );
  BUFX2 U16532 ( .A(n16089), .Y(n27183) );
  BUFX2 U16533 ( .A(n16168), .Y(n27184) );
  BUFX2 U16534 ( .A(n15938), .Y(n27185) );
  AND2X2 U16535 ( .A(n29478), .B(n25406), .Y(n34177) );
  INVX2 U16536 ( .A(n34177), .Y(n27186) );
  AND2X1 U16537 ( .A(n29652), .B(n34360), .Y(n16185) );
  INVX1 U16538 ( .A(n16185), .Y(n27187) );
  AND2X2 U16539 ( .A(n30040), .B(n29331), .Y(n32967) );
  INVX1 U16540 ( .A(n32967), .Y(n27188) );
  INVX2 U16541 ( .A(n32967), .Y(n27189) );
  AND2X2 U16542 ( .A(n29835), .B(n30002), .Y(n33792) );
  INVX1 U16543 ( .A(n33792), .Y(n27190) );
  INVX1 U16544 ( .A(n33792), .Y(n27191) );
  BUFX2 U16545 ( .A(n14675), .Y(n27192) );
  AND2X2 U16546 ( .A(n23611), .B(n34372), .Y(n16196) );
  INVX1 U16547 ( .A(n16196), .Y(n27193) );
  AND2X2 U16548 ( .A(n29807), .B(n32491), .Y(n33008) );
  INVX1 U16549 ( .A(n33008), .Y(n27194) );
  INVX1 U16550 ( .A(n33008), .Y(n27195) );
  BUFX2 U16551 ( .A(n30633), .Y(n27196) );
  AND2X2 U16552 ( .A(n27196), .B(n29207), .Y(n27300) );
  INVX1 U16553 ( .A(n27196), .Y(n34503) );
  AND2X2 U16554 ( .A(n30127), .B(T[0]), .Y(n34590) );
  INVX1 U16555 ( .A(n34590), .Y(n27197) );
  AND2X2 U16556 ( .A(n23299), .B(n32491), .Y(n33004) );
  INVX1 U16557 ( .A(n33004), .Y(n27198) );
  INVX1 U16558 ( .A(n33004), .Y(n27199) );
  INVX1 U16559 ( .A(n33004), .Y(n27200) );
  AND2X2 U16560 ( .A(n27248), .B(n27314), .Y(n29966) );
  INVX1 U16561 ( .A(n29966), .Y(n27201) );
  AND2X2 U16562 ( .A(n27248), .B(n27294), .Y(n29806) );
  INVX1 U16563 ( .A(n29806), .Y(n27202) );
  AND2X2 U16564 ( .A(n23289), .B(n21106), .Y(n33842) );
  INVX1 U16565 ( .A(n33842), .Y(n27203) );
  INVX1 U16566 ( .A(n33842), .Y(n27204) );
  INVX1 U16567 ( .A(n33842), .Y(n27205) );
  INVX1 U16568 ( .A(n33842), .Y(n27206) );
  AND2X2 U16569 ( .A(n27252), .B(n30626), .Y(n33661) );
  AND2X2 U16570 ( .A(n27294), .B(n21211), .Y(n27252) );
  INVX1 U16571 ( .A(n30027), .Y(n27208) );
  AND2X2 U16572 ( .A(n27213), .B(n27212), .Y(n8055) );
  INVX1 U16573 ( .A(n8055), .Y(n27209) );
  INVX2 U16574 ( .A(n8055), .Y(n27210) );
  INVX1 U16575 ( .A(n8055), .Y(n27211) );
  BUFX2 U16576 ( .A(n29500), .Y(n27212) );
  BUFX2 U16577 ( .A(n29501), .Y(n27213) );
  INVX2 U16578 ( .A(n29436), .Y(n29435) );
  INVX1 U16579 ( .A(n29319), .Y(n29315) );
  INVX2 U16580 ( .A(n2248), .Y(n28992) );
  INVX1 U16581 ( .A(n27152), .Y(n32101) );
  INVX1 U16582 ( .A(net106017), .Y(alt14_net96306) );
  INVX1 U16583 ( .A(net90071), .Y(alt14_net96326) );
  INVX8 U16584 ( .A(n29463), .Y(n29462) );
  INVX2 U16585 ( .A(n29393), .Y(n29387) );
  AND2X2 U16586 ( .A(n33056), .B(n33055), .Y(n27251) );
  AND2X2 U16587 ( .A(n25707), .B(n33052), .Y(n27255) );
  INVX1 U16588 ( .A(n31907), .Y(n29275) );
  INVX1 U16589 ( .A(n31908), .Y(n29276) );
  AND2X1 U16590 ( .A(n31868), .B(n29318), .Y(n27260) );
  AND2X1 U16591 ( .A(n27242), .B(n27304), .Y(n27262) );
  INVX1 U16592 ( .A(n30482), .Y(n29322) );
  INVX1 U16593 ( .A(n29248), .Y(n29243) );
  INVX1 U16594 ( .A(n29248), .Y(n27215) );
  INVX1 U16595 ( .A(n12071), .Y(n33203) );
  INVX1 U16596 ( .A(n12073), .Y(n33196) );
  INVX1 U16597 ( .A(n29468), .Y(n29467) );
  INVX1 U16598 ( .A(n25413), .Y(n29274) );
  INVX1 U16599 ( .A(n12067), .Y(n33226) );
  INVX1 U16600 ( .A(n12065), .Y(n33233) );
  INVX1 U16601 ( .A(n12049), .Y(n33318) );
  INVX1 U16602 ( .A(n12047), .Y(n33325) );
  INVX1 U16603 ( .A(n12043), .Y(n33349) );
  INVX1 U16604 ( .A(n12041), .Y(n33356) );
  INVX1 U16605 ( .A(n12037), .Y(n33379) );
  INVX1 U16606 ( .A(n12029), .Y(n33416) );
  INVX1 U16607 ( .A(n12061), .Y(n33257) );
  INVX1 U16608 ( .A(n12059), .Y(n33264) );
  INVX1 U16609 ( .A(n12055), .Y(n33287) );
  INVX1 U16610 ( .A(n12053), .Y(n33294) );
  INVX1 U16611 ( .A(n12035), .Y(n33386) );
  INVX1 U16612 ( .A(n12031), .Y(n33409) );
  INVX1 U16613 ( .A(n12077), .Y(n34346) );
  INVX1 U16614 ( .A(n34219), .Y(n29357) );
  INVX1 U16615 ( .A(n33885), .Y(n29346) );
  INVX1 U16616 ( .A(n34219), .Y(n29358) );
  INVX1 U16617 ( .A(n33885), .Y(n29347) );
  INVX1 U16618 ( .A(n29412), .Y(n29410) );
  INVX1 U16619 ( .A(n29403), .Y(n29401) );
  INVX1 U16620 ( .A(n29420), .Y(n29418) );
  INVX1 U16621 ( .A(n29452), .Y(n29451) );
  AND2X2 U16622 ( .A(oc[3]), .B(n29706), .Y(n27313) );
  INVX1 U16623 ( .A(n29252), .Y(n29251) );
  INVX1 U16624 ( .A(n29395), .Y(n29394) );
  INVX1 U16625 ( .A(n2253), .Y(n29465) );
  INVX1 U16626 ( .A(n29438), .Y(n29429) );
  INVX1 U16627 ( .A(n29439), .Y(n29425) );
  INVX1 U16628 ( .A(n29438), .Y(n29428) );
  INVX1 U16629 ( .A(n29437), .Y(n29430) );
  INVX1 U16630 ( .A(n29439), .Y(n29426) );
  INVX1 U16631 ( .A(n29438), .Y(n29427) );
  INVX1 U16632 ( .A(n29437), .Y(n29431) );
  INVX1 U16633 ( .A(n29437), .Y(n29432) );
  INVX1 U16634 ( .A(n29436), .Y(n29434) );
  INVX1 U16635 ( .A(n29436), .Y(n29433) );
  INVX1 U16636 ( .A(n29373), .Y(n29367) );
  INVX1 U16637 ( .A(n29373), .Y(n29368) );
  INVX1 U16638 ( .A(n29375), .Y(n29365) );
  INVX1 U16639 ( .A(alt14_net96268), .Y(alt14_net96250) );
  INVX1 U16640 ( .A(n25624), .Y(n27906) );
  INVX1 U16641 ( .A(n23191), .Y(n30841) );
  INVX1 U16642 ( .A(n23156), .Y(n30820) );
  INVX1 U16643 ( .A(n23157), .Y(n30860) );
  INVX1 U16644 ( .A(n34224), .Y(n29436) );
  INVX1 U16645 ( .A(n34224), .Y(n29437) );
  INVX1 U16646 ( .A(n34224), .Y(n29439) );
  INVX1 U16647 ( .A(n34224), .Y(n29438) );
  INVX1 U16648 ( .A(n29281), .Y(n29278) );
  INVX1 U16649 ( .A(n29281), .Y(n29279) );
  INVX1 U16650 ( .A(n29319), .Y(n29316) );
  INVX1 U16651 ( .A(n29319), .Y(n29317) );
  INVX1 U16652 ( .A(net96584), .Y(net96564) );
  INVX1 U16653 ( .A(net96584), .Y(net96566) );
  INVX1 U16654 ( .A(net96584), .Y(net96562) );
  INVX1 U16655 ( .A(net96582), .Y(net96570) );
  INVX1 U16656 ( .A(net96586), .Y(net96560) );
  INVX1 U16657 ( .A(net96582), .Y(net96568) );
  INVX1 U16658 ( .A(net96582), .Y(net96572) );
  INVX1 U16659 ( .A(n29385), .Y(n29373) );
  INVX1 U16660 ( .A(n29297), .Y(n29295) );
  INVX1 U16661 ( .A(n29297), .Y(n29294) );
  INVX1 U16662 ( .A(n29298), .Y(n29293) );
  INVX1 U16663 ( .A(n29298), .Y(n29292) );
  INVX1 U16664 ( .A(n29298), .Y(n29291) );
  INVX1 U16665 ( .A(n29384), .Y(n29375) );
  INVX1 U16666 ( .A(n29384), .Y(n29374) );
  INVX1 U16667 ( .A(n29281), .Y(n29280) );
  INVX1 U16668 ( .A(n29297), .Y(n29296) );
  INVX1 U16669 ( .A(alt14_net96258), .Y(alt14_net96268) );
  INVX1 U16670 ( .A(n28594), .Y(n28596) );
  INVX1 U16671 ( .A(n27906), .Y(n27905) );
  INVX1 U16672 ( .A(n21102), .Y(n28598) );
  INVX1 U16673 ( .A(alt14_net96306), .Y(alt14_net96304) );
  INVX1 U16674 ( .A(n28988), .Y(n28982) );
  INVX1 U16675 ( .A(n23149), .Y(n30721) );
  INVX1 U16676 ( .A(n23118), .Y(n30801) );
  INVX1 U16677 ( .A(n23136), .Y(n31388) );
  INVX1 U16678 ( .A(n23115), .Y(n31506) );
  INVX1 U16679 ( .A(n23127), .Y(n31586) );
  INVX1 U16680 ( .A(n23184), .Y(n31757) );
  INVX1 U16681 ( .A(n23129), .Y(n31797) );
  INVX1 U16682 ( .A(n23151), .Y(n30761) );
  INVX1 U16683 ( .A(n23171), .Y(n31429) );
  INVX1 U16684 ( .A(n23146), .Y(n30678) );
  INVX1 U16685 ( .A(n23148), .Y(n30701) );
  INVX1 U16686 ( .A(n23150), .Y(n30740) );
  INVX1 U16687 ( .A(n23154), .Y(n30780) );
  INVX1 U16688 ( .A(n23169), .Y(n31408) );
  INVX1 U16689 ( .A(n23161), .Y(n31057) );
  INVX1 U16690 ( .A(n23176), .Y(n31545) );
  INVX1 U16691 ( .A(n23180), .Y(n31680) );
  INVX1 U16692 ( .A(n23186), .Y(n31877) );
  INVX1 U16693 ( .A(n23159), .Y(n31019) );
  INVX1 U16694 ( .A(n23163), .Y(n31097) );
  INVX1 U16695 ( .A(n23175), .Y(n31525) );
  INVX1 U16696 ( .A(n23179), .Y(n31565) );
  INVX1 U16697 ( .A(n21487), .Y(n31605) );
  INVX1 U16698 ( .A(n23181), .Y(n31719) );
  INVX1 U16699 ( .A(n23034), .Y(n31275) );
  INVX1 U16700 ( .A(n23030), .Y(n31235) );
  INVX1 U16701 ( .A(n23027), .Y(n31195) );
  INVX1 U16702 ( .A(n23024), .Y(n31157) );
  INVX1 U16703 ( .A(n23017), .Y(n31039) );
  INVX1 U16704 ( .A(n23019), .Y(n31078) );
  INVX1 U16705 ( .A(n23022), .Y(n31118) );
  INVX1 U16706 ( .A(n23048), .Y(n31625) );
  INVX1 U16707 ( .A(n23058), .Y(n31739) );
  INVX1 U16708 ( .A(n23066), .Y(n31856) );
  INVX1 U16709 ( .A(n23055), .Y(n31700) );
  INVX1 U16710 ( .A(n23051), .Y(n31662) );
  INVX1 U16711 ( .A(n23060), .Y(n31778) );
  INVX1 U16712 ( .A(n23063), .Y(n31817) );
  INVX1 U16713 ( .A(n23076), .Y(n30664) );
  INVX1 U16714 ( .A(alt14_net96306), .Y(alt14_net96302) );
  INVX1 U16715 ( .A(n29195), .Y(n29230) );
  INVX1 U16716 ( .A(n28988), .Y(n28984) );
  INVX1 U16717 ( .A(n26181), .Y(n28985) );
  INVX1 U16718 ( .A(n26180), .Y(n28986) );
  INVX1 U16719 ( .A(n28988), .Y(n28983) );
  INVX1 U16720 ( .A(n26277), .Y(n29228) );
  INVX1 U16721 ( .A(n26715), .Y(n32235) );
  INVX1 U16722 ( .A(n26762), .Y(n32240) );
  INVX1 U16723 ( .A(n26936), .Y(n32245) );
  INVX1 U16724 ( .A(n26876), .Y(n32250) );
  INVX1 U16725 ( .A(n27093), .Y(n32265) );
  INVX1 U16726 ( .A(n27091), .Y(n32271) );
  INVX1 U16727 ( .A(n27221), .Y(n29298) );
  INVX1 U16728 ( .A(n27221), .Y(n29297) );
  INVX1 U16729 ( .A(n31862), .Y(n29281) );
  INVX1 U16730 ( .A(n31862), .Y(n29282) );
  INVX1 U16731 ( .A(n29305), .Y(n29302) );
  INVX1 U16732 ( .A(n29306), .Y(n29301) );
  INVX1 U16733 ( .A(n29306), .Y(n29300) );
  INVX1 U16734 ( .A(n29306), .Y(n29299) );
  INVX1 U16735 ( .A(n29305), .Y(n29303) );
  INVX1 U16736 ( .A(net96598), .Y(net96582) );
  INVX1 U16737 ( .A(net96600), .Y(net96586) );
  INVX1 U16738 ( .A(n29226), .Y(n29224) );
  INVX1 U16739 ( .A(net96598), .Y(net96592) );
  INVX1 U16740 ( .A(n29227), .Y(n29223) );
  INVX1 U16741 ( .A(n29227), .Y(n29222) );
  INVX1 U16742 ( .A(n29305), .Y(n29304) );
  INVX1 U16743 ( .A(n29226), .Y(n29225) );
  INVX1 U16744 ( .A(net96598), .Y(net96596) );
  INVX1 U16745 ( .A(n29442), .Y(n29440) );
  INVX1 U16746 ( .A(n29442), .Y(n29441) );
  INVX1 U16747 ( .A(n22967), .Y(n33076) );
  INVX1 U16748 ( .A(n25445), .Y(n32961) );
  INVX1 U16749 ( .A(n21222), .Y(n32777) );
  INVX1 U16750 ( .A(n27188), .Y(n32764) );
  INVX1 U16751 ( .A(n34420), .Y(n34417) );
  INVX1 U16752 ( .A(n25393), .Y(n32957) );
  INVX1 U16753 ( .A(n31894), .Y(n29195) );
  INVX1 U16754 ( .A(n28987), .Y(n28988) );
  INVX1 U16755 ( .A(n27224), .Y(n29313) );
  INVX1 U16756 ( .A(n29462), .Y(n28602) );
  INVX1 U16757 ( .A(n23189), .Y(n30690) );
  INVX1 U16758 ( .A(n23003), .Y(n30749) );
  INVX1 U16759 ( .A(n23005), .Y(n30789) );
  INVX1 U16760 ( .A(n23007), .Y(n30829) );
  INVX1 U16761 ( .A(n23192), .Y(n30869) );
  INVX1 U16762 ( .A(n23195), .Y(n31028) );
  INVX1 U16763 ( .A(n23018), .Y(n31066) );
  INVX1 U16764 ( .A(n23196), .Y(n31106) );
  INVX1 U16765 ( .A(n23041), .Y(n31438) );
  INVX1 U16766 ( .A(n23046), .Y(n31614) );
  INVX1 U16767 ( .A(n23040), .Y(n31417) );
  INVX1 U16768 ( .A(n25842), .Y(n31495) );
  INVX1 U16769 ( .A(n23045), .Y(n31554) );
  INVX1 U16770 ( .A(n23199), .Y(n31574) );
  INVX1 U16771 ( .A(n23049), .Y(n31650) );
  INVX1 U16772 ( .A(n22999), .Y(n31728) );
  INVX1 U16773 ( .A(n23013), .Y(n30971) );
  INVX1 U16774 ( .A(n23014), .Y(n30991) );
  INVX1 U16775 ( .A(n23023), .Y(n31146) );
  INVX1 U16776 ( .A(n23009), .Y(n30890) );
  INVX1 U16777 ( .A(n23010), .Y(n30910) );
  INVX1 U16778 ( .A(n23012), .Y(n30950) );
  INVX1 U16779 ( .A(n23025), .Y(n31183) );
  INVX1 U16780 ( .A(n23037), .Y(n31357) );
  INVX1 U16781 ( .A(n23028), .Y(n31223) );
  INVX1 U16782 ( .A(n23032), .Y(n31263) );
  INVX1 U16783 ( .A(n23039), .Y(n31397) );
  INVX1 U16784 ( .A(n23043), .Y(n31477) );
  INVX1 U16785 ( .A(n23059), .Y(n31766) );
  INVX1 U16786 ( .A(n29697), .Y(n32191) );
  INVX1 U16787 ( .A(n23020), .Y(n31125) );
  INVX1 U16788 ( .A(n26972), .Y(n31085) );
  INVX1 U16789 ( .A(n23062), .Y(n31824) );
  INVX1 U16790 ( .A(n26973), .Y(n31202) );
  INVX1 U16791 ( .A(n23029), .Y(n31242) );
  INVX1 U16792 ( .A(n26971), .Y(n31785) );
  INVX1 U16793 ( .A(n23054), .Y(n31707) );
  INVX1 U16794 ( .A(n25768), .Y(n33082) );
  INVX1 U16795 ( .A(n26304), .Y(n28603) );
  INVX1 U16796 ( .A(n27224), .Y(n29314) );
  INVX1 U16797 ( .A(n25624), .Y(n27903) );
  INVX1 U16798 ( .A(n29464), .Y(n28601) );
  INVX1 U16799 ( .A(n29464), .Y(n28600) );
  INVX1 U16800 ( .A(n25448), .Y(n32463) );
  AND2X1 U16801 ( .A(n27242), .B(n23443), .Y(n27221) );
  INVX1 U16802 ( .A(n27106), .Y(n32438) );
  INVX1 U16803 ( .A(n26943), .Y(n32446) );
  INVX1 U16804 ( .A(n27109), .Y(n32319) );
  INVX1 U16805 ( .A(n27009), .Y(n32415) );
  INVX1 U16806 ( .A(n27112), .Y(n32295) );
  INVX1 U16807 ( .A(n27012), .Y(n32327) );
  INVX1 U16808 ( .A(n26944), .Y(n32423) );
  INVX1 U16809 ( .A(n26947), .Y(n32335) );
  INVX1 U16810 ( .A(n27015), .Y(n32303) );
  BUFX2 U16811 ( .A(n27147), .Y(n29211) );
  INVX1 U16812 ( .A(n25398), .Y(n34495) );
  INVX1 U16813 ( .A(n26934), .Y(n32200) );
  INVX1 U16814 ( .A(n27089), .Y(n32205) );
  INVX1 U16815 ( .A(n26815), .Y(n32210) );
  INVX1 U16816 ( .A(n27003), .Y(n32255) );
  INVX1 U16817 ( .A(n26817), .Y(n32260) );
  INVX1 U16818 ( .A(n27087), .Y(n32215) );
  INVX1 U16819 ( .A(n26760), .Y(n32220) );
  INVX1 U16820 ( .A(n26872), .Y(n32279) );
  INVX1 U16821 ( .A(n26813), .Y(n32311) );
  INVX1 U16822 ( .A(n25382), .Y(n32407) );
  INVX1 U16823 ( .A(n27001), .Y(n32225) );
  INVX1 U16824 ( .A(n26874), .Y(n32230) );
  INVX1 U16825 ( .A(n26758), .Y(n32287) );
  INVX1 U16826 ( .A(n25434), .Y(n34496) );
  INVX1 U16827 ( .A(n25283), .Y(n32363) );
  INVX1 U16828 ( .A(n25308), .Y(n32427) );
  INVX1 U16829 ( .A(n25269), .Y(n32331) );
  INVX1 U16830 ( .A(n25273), .Y(n32343) );
  INVX1 U16831 ( .A(n25277), .Y(n32351) );
  INVX1 U16832 ( .A(n25236), .Y(n32224) );
  INVX1 U16833 ( .A(n25226), .Y(n32199) );
  INVX1 U16834 ( .A(n25230), .Y(n32209) );
  INVX1 U16835 ( .A(n25238), .Y(n32229) );
  INVX1 U16836 ( .A(n25315), .Y(n32457) );
  INVX1 U16837 ( .A(n25309), .Y(n32434) );
  INVX1 U16838 ( .A(n25271), .Y(n32339) );
  INVX1 U16839 ( .A(n25302), .Y(n32403) );
  INVX1 U16840 ( .A(n25263), .Y(n32307) );
  INVX1 U16841 ( .A(n25285), .Y(n32367) );
  INVX1 U16842 ( .A(n27234), .Y(n29306) );
  INVX1 U16843 ( .A(n27234), .Y(n29305) );
  INVX1 U16844 ( .A(n27235), .Y(n29226) );
  INVX1 U16845 ( .A(alt5_net95670), .Y(alt5_net95656) );
  INVX1 U16846 ( .A(alt5_net95668), .Y(alt5_net95652) );
  INVX1 U16847 ( .A(n27235), .Y(n29227) );
  INVX1 U16848 ( .A(n29290), .Y(n29285) );
  INVX1 U16849 ( .A(n29290), .Y(n29283) );
  INVX1 U16850 ( .A(n29290), .Y(n29284) );
  INVX1 U16851 ( .A(n29289), .Y(n29286) );
  INVX1 U16852 ( .A(n29312), .Y(n29310) );
  INVX1 U16853 ( .A(n29312), .Y(n29309) );
  INVX1 U16854 ( .A(n29312), .Y(n29307) );
  INVX1 U16855 ( .A(n29312), .Y(n29308) );
  INVX1 U16856 ( .A(n29289), .Y(n29288) );
  INVX1 U16857 ( .A(n29312), .Y(n29311) );
  INVX1 U16858 ( .A(net96604), .Y(net96600) );
  INVX1 U16859 ( .A(net96604), .Y(net96598) );
  INVX1 U16860 ( .A(n31892), .Y(n29255) );
  INVX1 U16861 ( .A(n31892), .Y(n29257) );
  INVX1 U16862 ( .A(n31892), .Y(n29258) );
  INVX1 U16863 ( .A(n31892), .Y(n29256) );
  INVX1 U16864 ( .A(n31892), .Y(n29254) );
  INVX1 U16865 ( .A(n27271), .Y(n29260) );
  INVX1 U16866 ( .A(n27271), .Y(n29262) );
  INVX1 U16867 ( .A(n27271), .Y(n29263) );
  INVX1 U16868 ( .A(n29265), .Y(n29264) );
  INVX1 U16869 ( .A(n29241), .Y(n29240) );
  INVX1 U16870 ( .A(n29460), .Y(n29453) );
  INVX1 U16871 ( .A(n29460), .Y(n29454) );
  INVX1 U16872 ( .A(n29460), .Y(n29455) );
  INVX1 U16873 ( .A(n29459), .Y(n29456) );
  INVX1 U16874 ( .A(n29459), .Y(n29457) );
  INVX1 U16875 ( .A(n29459), .Y(n29458) );
  INVX1 U16876 ( .A(n31892), .Y(n29259) );
  INVX1 U16877 ( .A(n29471), .Y(n27700) );
  INVX1 U16878 ( .A(n29471), .Y(n27701) );
  INVX1 U16879 ( .A(n34263), .Y(n34273) );
  INVX1 U16880 ( .A(n25317), .Y(n34260) );
  AND2X2 U16881 ( .A(n27019), .B(net114546), .Y(n27223) );
  AND2X2 U16882 ( .A(n20995), .B(n27152), .Y(n27224) );
  INVX1 U16883 ( .A(n34407), .Y(n34414) );
  INVX1 U16884 ( .A(n34334), .Y(n34332) );
  INVX1 U16885 ( .A(net53601), .Y(alt14_net55935) );
  INVX1 U16886 ( .A(net53601), .Y(alt14_net55927) );
  INVX1 U16887 ( .A(net53601), .Y(alt14_net55921) );
  INVX1 U16888 ( .A(n22972), .Y(n34264) );
  INVX1 U16889 ( .A(n34326), .Y(n34410) );
  AND2X1 U16890 ( .A(n31618), .B(net96340), .Y(n27226) );
  AND2X1 U16891 ( .A(n31732), .B(net96340), .Y(n27227) );
  AND2X1 U16892 ( .A(n31150), .B(net96340), .Y(n27228) );
  AND2X1 U16893 ( .A(n31848), .B(net96340), .Y(n27229) );
  AND2X1 U16894 ( .A(n30995), .B(net96340), .Y(n27230) );
  AND2X1 U16895 ( .A(n31032), .B(net96340), .Y(n27231) );
  XNOR2X1 U16896 ( .A(n26053), .B(n29206), .Y(n27233) );
  INVX1 U16897 ( .A(n22964), .Y(n28991) );
  INVX1 U16898 ( .A(n25644), .Y(n34319) );
  INVX1 U16899 ( .A(n34418), .Y(n34421) );
  INVX1 U16900 ( .A(n29467), .Y(n28990) );
  INVX1 U16901 ( .A(n25455), .Y(n33531) );
  INVX1 U16902 ( .A(n27026), .Y(n33748) );
  INVX1 U16903 ( .A(n27206), .Y(n33861) );
  INVX1 U16904 ( .A(n27120), .Y(n33815) );
  INVX1 U16905 ( .A(n21384), .Y(n33417) );
  INVX1 U16906 ( .A(n21387), .Y(n33234) );
  AND2X1 U16907 ( .A(n27247), .B(n29352), .Y(n27234) );
  AND2X1 U16908 ( .A(n30482), .B(net96340), .Y(n27235) );
  BUFX2 U16909 ( .A(n25621), .Y(n27916) );
  INVX1 U16910 ( .A(n30111), .Y(n30451) );
  INVX1 U16911 ( .A(n21378), .Y(n33784) );
  BUFX2 U16912 ( .A(n27146), .Y(n29210) );
  INVX1 U16913 ( .A(n25279), .Y(n32355) );
  INVX1 U16914 ( .A(n25281), .Y(n32359) );
  INVX1 U16915 ( .A(n25294), .Y(n32387) );
  INVX1 U16916 ( .A(n25298), .Y(n32395) );
  INVX1 U16917 ( .A(n25296), .Y(n32391) );
  INVX1 U16918 ( .A(n25252), .Y(n32264) );
  INVX1 U16919 ( .A(n25250), .Y(n32259) );
  INVX1 U16920 ( .A(n25248), .Y(n32254) );
  INVX1 U16921 ( .A(n25306), .Y(n32419) );
  INVX1 U16922 ( .A(n25267), .Y(n32323) );
  INVX1 U16923 ( .A(n25260), .Y(n32291) );
  INVX1 U16924 ( .A(n25261), .Y(n32299) );
  INVX1 U16925 ( .A(n25289), .Y(n32375) );
  INVX1 U16926 ( .A(n25242), .Y(n32239) );
  INVX1 U16927 ( .A(n25275), .Y(n32347) );
  INVX1 U16928 ( .A(n25290), .Y(n32379) );
  INVX1 U16929 ( .A(n25244), .Y(n32244) );
  INVX1 U16930 ( .A(n25304), .Y(n32411) );
  INVX1 U16931 ( .A(n25265), .Y(n32315) );
  INVX1 U16932 ( .A(n25258), .Y(n32283) );
  INVX1 U16933 ( .A(n25292), .Y(n32383) );
  INVX1 U16934 ( .A(n25246), .Y(n32249) );
  INVX1 U16935 ( .A(n25228), .Y(n32204) );
  INVX1 U16936 ( .A(n25232), .Y(n32214) );
  INVX1 U16937 ( .A(n25234), .Y(n32219) );
  INVX1 U16938 ( .A(n25313), .Y(n32450) );
  INVX1 U16939 ( .A(n25311), .Y(n32442) );
  INVX1 U16940 ( .A(n25287), .Y(n32371) );
  INVX1 U16941 ( .A(n25240), .Y(n32234) );
  INVX1 U16942 ( .A(n25256), .Y(n32275) );
  INVX1 U16943 ( .A(n25300), .Y(n32399) );
  INVX1 U16944 ( .A(n25254), .Y(n32270) );
  INVX1 U16945 ( .A(n30136), .Y(n30476) );
  INVX1 U16946 ( .A(n30102), .Y(n30442) );
  INVX1 U16947 ( .A(n30093), .Y(n30433) );
  INVX1 U16948 ( .A(n30128), .Y(n30464) );
  AND2X2 U16949 ( .A(n27244), .B(net147379), .Y(n27240) );
  INVX1 U16950 ( .A(n27259), .Y(n29460) );
  INVX1 U16951 ( .A(n27259), .Y(n29459) );
  INVX1 U16952 ( .A(n27260), .Y(n29289) );
  INVX1 U16953 ( .A(n27260), .Y(n29290) );
  INVX1 U16954 ( .A(n27261), .Y(n29270) );
  INVX1 U16955 ( .A(n26051), .Y(n29184) );
  INVX1 U16956 ( .A(n27261), .Y(n29271) );
  AND2X2 U16957 ( .A(n25211), .B(net96340), .Y(net102091) );
  INVX1 U16958 ( .A(n27271), .Y(n29265) );
  AND2X1 U16959 ( .A(n31914), .B(n29381), .Y(n27242) );
  AND2X1 U16960 ( .A(n33995), .B(n33996), .Y(n27245) );
  AND2X1 U16961 ( .A(net53623), .B(net53601), .Y(n27246) );
  INVX1 U16962 ( .A(n29242), .Y(n29237) );
  INVX1 U16963 ( .A(n21438), .Y(n29242) );
  INVX1 U16964 ( .A(n29242), .Y(n29239) );
  INVX1 U16965 ( .A(n29242), .Y(n29238) );
  INVX1 U16966 ( .A(n21438), .Y(n29241) );
  INVX1 U16967 ( .A(n29322), .Y(n29321) );
  INVX1 U16968 ( .A(n29452), .Y(n29444) );
  INVX1 U16969 ( .A(n29452), .Y(n29445) );
  INVX1 U16970 ( .A(n29452), .Y(n29446) );
  INVX1 U16971 ( .A(n29450), .Y(n29447) );
  INVX1 U16972 ( .A(n29450), .Y(n29448) );
  INVX1 U16973 ( .A(n29450), .Y(n29449) );
  AND2X1 U16974 ( .A(n31914), .B(net96340), .Y(n27247) );
  INVX1 U16975 ( .A(n15921), .Y(n34506) );
  INVX1 U16976 ( .A(n15931), .Y(n34589) );
  INVX1 U16977 ( .A(n15923), .Y(n34586) );
  INVX1 U16978 ( .A(n26868), .Y(n34576) );
  INVX1 U16979 ( .A(n25219), .Y(n34596) );
  INVX1 U16980 ( .A(n26970), .Y(n30087) );
  INVX1 U16981 ( .A(n26672), .Y(n30149) );
  INVX1 U16982 ( .A(n26784), .Y(n30289) );
  INVX1 U16983 ( .A(n26845), .Y(n30104) );
  INVX1 U16984 ( .A(n26742), .Y(n30121) );
  INVX1 U16985 ( .A(n26673), .Y(n30138) );
  INVX1 U16986 ( .A(n26617), .Y(n30159) );
  INVX1 U16987 ( .A(n26592), .Y(n30169) );
  INVX1 U16988 ( .A(n26844), .Y(n30180) );
  INVX1 U16989 ( .A(n26702), .Y(n30299) );
  INVX1 U16990 ( .A(n26641), .Y(n30309) );
  INVX1 U16991 ( .A(n26967), .Y(n30322) );
  INVX1 U16992 ( .A(n27052), .Y(n30195) );
  INVX1 U16993 ( .A(n26786), .Y(n30205) );
  INVX1 U16994 ( .A(n26703), .Y(n30215) );
  INVX1 U16995 ( .A(n26904), .Y(n30229) );
  INVX1 U16996 ( .A(n33555), .Y(n29882) );
  INVX1 U16997 ( .A(n30557), .Y(n29897) );
  INVX1 U16998 ( .A(n27715), .Y(n27711) );
  INVX1 U16999 ( .A(n27715), .Y(n27710) );
  INVX1 U17000 ( .A(n27715), .Y(n27714) );
  INVX1 U17001 ( .A(n27715), .Y(n27713) );
  INVX1 U17002 ( .A(n27715), .Y(n27712) );
  INVX1 U17003 ( .A(n27715), .Y(n27706) );
  INVX1 U17004 ( .A(n27715), .Y(n27705) );
  INVX1 U17005 ( .A(n27715), .Y(n27709) );
  INVX1 U17006 ( .A(n27715), .Y(n27708) );
  INVX1 U17007 ( .A(n27715), .Y(n27707) );
  INVX1 U17008 ( .A(n27703), .Y(n27704) );
  INVX1 U17009 ( .A(n22990), .Y(n30076) );
  INVX1 U17010 ( .A(n27062), .Y(n29320) );
  INVX1 U17011 ( .A(n29700), .Y(n34555) );
  INVX1 U17012 ( .A(n29885), .Y(n29894) );
  INVX1 U17013 ( .A(n29218), .Y(n29217) );
  INVX1 U17014 ( .A(n30485), .Y(n29633) );
  INVX1 U17015 ( .A(n25395), .Y(n33120) );
  INVX2 U17016 ( .A(n26269), .Y(n33277) );
  INVX1 U17017 ( .A(n30066), .Y(n30046) );
  INVX1 U17018 ( .A(n13803), .Y(n29624) );
  INVX1 U17019 ( .A(n34423), .Y(n34424) );
  INVX1 U17020 ( .A(n25420), .Y(n30410) );
  BUFX2 U17021 ( .A(n25450), .Y(n28609) );
  BUFX2 U17022 ( .A(n25450), .Y(n28608) );
  BUFX2 U17023 ( .A(n2249), .Y(n28994) );
  INVX1 U17024 ( .A(n33163), .Y(n33161) );
  INVX1 U17025 ( .A(n25833), .Y(n34427) );
  INVX1 U17026 ( .A(net112859), .Y(net94645) );
  INVX1 U17027 ( .A(n22994), .Y(n29511) );
  INVX1 U17028 ( .A(net143010), .Y(net94647) );
  INVX1 U17029 ( .A(n34425), .Y(n34399) );
  INVX1 U17030 ( .A(n33140), .Y(n33148) );
  INVX1 U17031 ( .A(n25401), .Y(n33166) );
  AND2X2 U17032 ( .A(n21556), .B(n26788), .Y(n27253) );
  INVX1 U17033 ( .A(n33091), .Y(n33087) );
  INVX1 U17034 ( .A(n33106), .Y(n33146) );
  INVX1 U17035 ( .A(n33097), .Y(n33095) );
  INVX1 U17036 ( .A(n25071), .Y(n33086) );
  INVX1 U17037 ( .A(n24985), .Y(n33110) );
  INVX1 U17038 ( .A(n22993), .Y(n34365) );
  INVX1 U17039 ( .A(n33071), .Y(n33092) );
  INVX1 U17040 ( .A(n22983), .Y(n34198) );
  INVX1 U17041 ( .A(n22995), .Y(n34199) );
  INVX1 U17042 ( .A(n34437), .Y(n34231) );
  INVX1 U17043 ( .A(n8036), .Y(n30044) );
  XNOR2X1 U17044 ( .A(n25420), .B(n21186), .Y(n27254) );
  MUX2X1 U17045 ( .B(n28039), .A(n28038), .S(net53623), .Y(n4227) );
  INVX1 U17046 ( .A(n29247), .Y(n29244) );
  INVX1 U17047 ( .A(n29247), .Y(n29245) );
  INVX1 U17048 ( .A(n29247), .Y(n29246) );
  INVX1 U17049 ( .A(n29274), .Y(n29272) );
  INVX1 U17050 ( .A(n29274), .Y(n29273) );
  INVX1 U17051 ( .A(n29467), .Y(n28989) );
  INVX1 U17052 ( .A(n27211), .Y(n33996) );
  INVX1 U17053 ( .A(n27200), .Y(n34342) );
  INVX1 U17054 ( .A(n25450), .Y(n33995) );
  AND2X1 U17055 ( .A(n34174), .B(net90055), .Y(n27259) );
  INVX1 U17056 ( .A(n30094), .Y(n30434) );
  INVX1 U17057 ( .A(n30129), .Y(n30465) );
  AND2X1 U17058 ( .A(n30086), .B(n34189), .Y(n27268) );
  INVX1 U17059 ( .A(n30283), .Y(n30321) );
  INVX1 U17060 ( .A(n30189), .Y(n30228) );
  AND2X1 U17061 ( .A(n27301), .B(n30127), .Y(n27269) );
  INVX1 U17062 ( .A(n30373), .Y(n30411) );
  INVX1 U17063 ( .A(n30328), .Y(n30364) );
  INVX1 U17064 ( .A(n30282), .Y(n30320) );
  INVX1 U17065 ( .A(n30236), .Y(n30273) );
  INVX1 U17066 ( .A(n30188), .Y(n30227) );
  INVX1 U17067 ( .A(n30329), .Y(n30365) );
  INVX1 U17068 ( .A(n30237), .Y(n30274) );
  INVX1 U17069 ( .A(n30119), .Y(n30458) );
  INVX1 U17070 ( .A(n30110), .Y(n30450) );
  INVX1 U17071 ( .A(n30374), .Y(n30412) );
  INVX1 U17072 ( .A(n30420), .Y(n30472) );
  INVX1 U17073 ( .A(n30419), .Y(n30475) );
  INVX1 U17074 ( .A(n21556), .Y(n29748) );
  INVX1 U17075 ( .A(n13801), .Y(n34170) );
  INVX1 U17076 ( .A(n21429), .Y(n34172) );
  INVX1 U17077 ( .A(n29178), .Y(n29183) );
  INVX1 U17078 ( .A(n2252), .Y(n29178) );
  INVX1 U17079 ( .A(n29346), .Y(n29344) );
  INVX1 U17080 ( .A(n29346), .Y(n29345) );
  INVX1 U17081 ( .A(n29357), .Y(n29356) );
  INVX1 U17082 ( .A(n29358), .Y(n29354) );
  INVX1 U17083 ( .A(n29413), .Y(n29406) );
  INVX1 U17084 ( .A(n29451), .Y(n29450) );
  INVX1 U17085 ( .A(n2251), .Y(alt5_net95676) );
  INVX1 U17086 ( .A(n29392), .Y(n29391) );
  INVX1 U17087 ( .A(n29216), .Y(n29214) );
  INVX1 U17088 ( .A(n29418), .Y(n29417) );
  INVX1 U17089 ( .A(reset), .Y(net96340) );
  INVX1 U17090 ( .A(n31868), .Y(n29221) );
  INVX1 U17091 ( .A(n16232), .Y(n34588) );
  INVX1 U17092 ( .A(n15948), .Y(n34570) );
  INVX1 U17093 ( .A(n16022), .Y(n34565) );
  INVX1 U17094 ( .A(n16099), .Y(n34580) );
  INVX1 U17095 ( .A(n16180), .Y(n34559) );
  INVX1 U17096 ( .A(n15989), .Y(n34577) );
  INVX1 U17097 ( .A(n16221), .Y(n34593) );
  INVX1 U17098 ( .A(n16195), .Y(n34502) );
  INVX1 U17099 ( .A(n27273), .Y(n30556) );
  INVX1 U17100 ( .A(n29653), .Y(n29654) );
  INVX1 U17101 ( .A(n16034), .Y(n34564) );
  INVX1 U17102 ( .A(n16192), .Y(n34558) );
  INVX1 U17103 ( .A(n15960), .Y(n34569) );
  INVX1 U17104 ( .A(n16111), .Y(n34579) );
  INVX1 U17105 ( .A(n29649), .Y(n34501) );
  INVX1 U17106 ( .A(n15963), .Y(n34499) );
  INVX1 U17107 ( .A(n16114), .Y(n34500) );
  INVX1 U17108 ( .A(n24979), .Y(n30051) );
  INVX1 U17109 ( .A(n16080), .Y(n34581) );
  INVX1 U17110 ( .A(n16154), .Y(n34560) );
  INVX1 U17111 ( .A(n15927), .Y(n34571) );
  INVX1 U17112 ( .A(n16003), .Y(n34566) );
  INVX1 U17113 ( .A(n16152), .Y(n34557) );
  INVX1 U17114 ( .A(n15925), .Y(n34568) );
  INVX1 U17115 ( .A(n16001), .Y(n34563) );
  INVX1 U17116 ( .A(n16078), .Y(n34578) );
  INVX1 U17117 ( .A(n26919), .Y(n34561) );
  INVX1 U17118 ( .A(n26859), .Y(n34567) );
  INVX1 U17119 ( .A(n27053), .Y(n30144) );
  INVX1 U17120 ( .A(n26969), .Y(n30190) );
  INVX1 U17121 ( .A(n26642), .Y(n30238) );
  INVX1 U17122 ( .A(n26842), .Y(n30284) );
  INVX1 U17123 ( .A(n26615), .Y(n30330) );
  INVX1 U17124 ( .A(n26590), .Y(n30335) );
  INVX1 U17125 ( .A(n26739), .Y(n30375) );
  INVX1 U17126 ( .A(n26906), .Y(n30095) );
  INVX1 U17127 ( .A(n26787), .Y(n30112) );
  INVX1 U17128 ( .A(n26704), .Y(n30130) );
  INVX1 U17129 ( .A(n26643), .Y(n30154) );
  INVX1 U17130 ( .A(n27150), .Y(n30164) );
  INVX1 U17131 ( .A(n26905), .Y(n30174) );
  INVX1 U17132 ( .A(n26843), .Y(n30200) );
  INVX1 U17133 ( .A(n26741), .Y(n30210) );
  INVX1 U17134 ( .A(n26671), .Y(n30220) );
  INVX1 U17135 ( .A(n27051), .Y(n30248) );
  INVX1 U17136 ( .A(n26968), .Y(n30258) );
  INVX1 U17137 ( .A(n26740), .Y(n30294) );
  INVX1 U17138 ( .A(n26670), .Y(n30304) );
  INVX1 U17139 ( .A(n27050), .Y(n30314) );
  INVX1 U17140 ( .A(n26966), .Y(n30340) );
  INVX1 U17141 ( .A(n26902), .Y(n30349) );
  INVX1 U17142 ( .A(n26841), .Y(n30354) );
  INVX1 U17143 ( .A(n26783), .Y(n30359) );
  INVX1 U17144 ( .A(n27049), .Y(n30366) );
  INVX1 U17145 ( .A(n26701), .Y(n30394) );
  INVX1 U17146 ( .A(n26640), .Y(n30404) );
  INVX1 U17147 ( .A(n26700), .Y(n30421) );
  INVX1 U17148 ( .A(n27148), .Y(n30435) );
  INVX1 U17149 ( .A(n26613), .Y(n30452) );
  INVX1 U17150 ( .A(n26588), .Y(n30466) );
  INVX1 U17151 ( .A(n26616), .Y(n30243) );
  INVX1 U17152 ( .A(n27149), .Y(n30380) );
  INVX1 U17153 ( .A(n26591), .Y(n30253) );
  INVX1 U17154 ( .A(n26903), .Y(n30263) );
  INVX1 U17155 ( .A(n26785), .Y(n30275) );
  INVX1 U17156 ( .A(n26669), .Y(n30389) );
  INVX1 U17157 ( .A(n26614), .Y(n30399) );
  INVX1 U17158 ( .A(n26589), .Y(n30413) );
  INVX1 U17159 ( .A(n26738), .Y(n30427) );
  INVX1 U17160 ( .A(n26639), .Y(n30444) );
  INVX1 U17161 ( .A(n27151), .Y(n30080) );
  INVX1 U17162 ( .A(n16066), .Y(n34595) );
  INVX1 U17163 ( .A(n16224), .Y(n34592) );
  INVX1 U17164 ( .A(n15992), .Y(n34575) );
  INVX1 U17165 ( .A(n16143), .Y(n34585) );
  INVX1 U17166 ( .A(n24932), .Y(n34606) );
  INVX1 U17167 ( .A(n24933), .Y(n34609) );
  INVX1 U17168 ( .A(n24934), .Y(n34599) );
  INVX1 U17169 ( .A(n24935), .Y(n34602) );
  INVX1 U17170 ( .A(n29470), .Y(n27702) );
  INVX1 U17171 ( .A(n24963), .Y(n34603) );
  INVX1 U17172 ( .A(n29328), .Y(n29325) );
  INVX1 U17173 ( .A(n29328), .Y(n29326) );
  INVX1 U17174 ( .A(n29329), .Y(n29323) );
  INVX1 U17175 ( .A(n29329), .Y(n29324) );
  INVX1 U17176 ( .A(n29729), .Y(n29738) );
  INVX1 U17177 ( .A(n29328), .Y(n29327) );
  AND2X1 U17178 ( .A(n29352), .B(n30550), .Y(n27275) );
  INVX1 U17179 ( .A(n29335), .Y(n29333) );
  INVX1 U17180 ( .A(n29335), .Y(n29332) );
  INVX1 U17181 ( .A(n20978), .Y(n27715) );
  INVX1 U17182 ( .A(n29335), .Y(n29334) );
  INVX1 U17183 ( .A(address[3]), .Y(n27703) );
  INVX1 U17184 ( .A(n33994), .Y(n22637) );
  INVX1 U17185 ( .A(n33932), .Y(n22626) );
  INVX1 U17186 ( .A(n33916), .Y(n22627) );
  INVX1 U17187 ( .A(n23096), .Y(n33114) );
  INVX1 U17188 ( .A(n25212), .Y(n30644) );
  AND2X2 U17189 ( .A(n30632), .B(n30631), .Y(n27276) );
  INVX1 U17190 ( .A(n33395), .Y(n33397) );
  INVX1 U17191 ( .A(n12033), .Y(n33396) );
  INVX1 U17192 ( .A(n33404), .Y(n33406) );
  INVX1 U17193 ( .A(n12032), .Y(n33405) );
  INVX1 U17194 ( .A(n33221), .Y(n33223) );
  INVX1 U17195 ( .A(n12068), .Y(n33222) );
  INVX1 U17196 ( .A(n33365), .Y(n33367) );
  INVX1 U17197 ( .A(n12039), .Y(n33366) );
  INVX1 U17198 ( .A(n33374), .Y(n33376) );
  INVX1 U17199 ( .A(n12038), .Y(n33375) );
  INVX1 U17200 ( .A(n33186), .Y(n33188) );
  INVX1 U17201 ( .A(n12074), .Y(n33187) );
  INVX1 U17202 ( .A(n33212), .Y(n33214) );
  INVX1 U17203 ( .A(n12069), .Y(n33213) );
  INVX1 U17204 ( .A(n34226), .Y(n34228) );
  INVX1 U17205 ( .A(n12075), .Y(n34227) );
  INVX1 U17206 ( .A(n33273), .Y(n33275) );
  INVX1 U17207 ( .A(n12057), .Y(n33274) );
  INVX1 U17208 ( .A(n33282), .Y(n33284) );
  INVX1 U17209 ( .A(n12056), .Y(n33283) );
  INVX1 U17210 ( .A(n33313), .Y(n33315) );
  INVX1 U17211 ( .A(n12050), .Y(n33314) );
  INVX1 U17212 ( .A(n33344), .Y(n33346) );
  INVX1 U17213 ( .A(n12044), .Y(n33345) );
  INVX1 U17214 ( .A(n33426), .Y(n33428) );
  INVX1 U17215 ( .A(n12027), .Y(n33427) );
  INVX1 U17216 ( .A(n33252), .Y(n33254) );
  INVX1 U17217 ( .A(n12062), .Y(n33253) );
  INVX1 U17218 ( .A(n33304), .Y(n33306) );
  INVX1 U17219 ( .A(n12051), .Y(n33305) );
  INVX1 U17220 ( .A(n33335), .Y(n33337) );
  INVX1 U17221 ( .A(n12045), .Y(n33336) );
  INVX1 U17222 ( .A(n33243), .Y(n33245) );
  INVX1 U17223 ( .A(n12063), .Y(n33244) );
  INVX1 U17224 ( .A(n25336), .Y(n33129) );
  AND2X2 U17225 ( .A(n29723), .B(n29706), .Y(n27294) );
  INVX1 U17226 ( .A(n23200), .Y(n29628) );
  INVX1 U17227 ( .A(n22985), .Y(n30685) );
  INVX1 U17228 ( .A(n25334), .Y(n29629) );
  INVX1 U17229 ( .A(n25406), .Y(n29510) );
  AND2X1 U17230 ( .A(n25331), .B(n25407), .Y(n27297) );
  INVX1 U17231 ( .A(n33918), .Y(n34209) );
  INVX1 U17232 ( .A(n25330), .Y(n29509) );
  INVX1 U17233 ( .A(n19664), .Y(n33919) );
  INVX1 U17234 ( .A(n19663), .Y(n33920) );
  INVX1 U17235 ( .A(n19662), .Y(n33917) );
  INVX1 U17236 ( .A(n23088), .Y(n29845) );
  INVX1 U17237 ( .A(n33133), .Y(n33131) );
  INVX1 U17238 ( .A(n25416), .Y(n34358) );
  INVX1 U17239 ( .A(n32892), .Y(n33052) );
  INVX1 U17240 ( .A(n32515), .Y(n33056) );
  INVX1 U17241 ( .A(n22966), .Y(n33051) );
  INVX1 U17242 ( .A(n32565), .Y(n33055) );
  AND2X1 U17243 ( .A(n32561), .B(n32560), .Y(n32562) );
  INVX1 U17244 ( .A(n24926), .Y(n30653) );
  INVX1 U17245 ( .A(n29251), .Y(n29249) );
  INVX1 U17246 ( .A(n29251), .Y(n29250) );
  AND2X2 U17247 ( .A(net103869), .B(n34338), .Y(n27304) );
  AND2X1 U17248 ( .A(n30086), .B(n23441), .Y(n27308) );
  INVX1 U17249 ( .A(n30187), .Y(n30226) );
  INVX1 U17250 ( .A(net103869), .Y(net90055) );
  INVX1 U17251 ( .A(n27172), .Y(n34612) );
  AND2X1 U17252 ( .A(n9146), .B(n29381), .Y(n21804) );
  AND2X1 U17253 ( .A(n9150), .B(n29381), .Y(n21808) );
  AND2X1 U17254 ( .A(n9156), .B(n29381), .Y(n21814) );
  INVX1 U17255 ( .A(n29188), .Y(n29186) );
  INVX1 U17256 ( .A(n29188), .Y(n29187) );
  INVX1 U17257 ( .A(n29420), .Y(n29419) );
  INVX1 U17258 ( .A(n22058), .Y(n29452) );
  INVX1 U17259 ( .A(n29403), .Y(n29402) );
  INVX1 U17260 ( .A(n29411), .Y(n29405) );
  INVX1 U17261 ( .A(n29412), .Y(n29411) );
  INVX1 U17262 ( .A(n29394), .Y(n29393) );
  INVX1 U17263 ( .A(n29394), .Y(n29392) );
  AND2X1 U17264 ( .A(n15177), .B(n30126), .Y(n27311) );
  AND2X1 U17265 ( .A(n30327), .B(n15174), .Y(n27312) );
  INVX1 U17266 ( .A(n30071), .Y(n30135) );
  INVX1 U17267 ( .A(n30072), .Y(n30418) );
  INVX1 U17268 ( .A(n15201), .Y(n33562) );
  INVX1 U17269 ( .A(n33561), .Y(n33563) );
  INVX1 U17270 ( .A(n27118), .Y(n34504) );
  INVX1 U17271 ( .A(n15169), .Y(n34598) );
  INVX1 U17272 ( .A(n15066), .Y(n34601) );
  INVX1 U17273 ( .A(n14968), .Y(n34605) );
  INVX1 U17274 ( .A(n14772), .Y(n34608) );
  INVX1 U17275 ( .A(n15998), .Y(n34562) );
  INVX1 U17276 ( .A(n15204), .Y(n34497) );
  INVX1 U17277 ( .A(n14348), .Y(n33992) );
  INVX1 U17278 ( .A(n32462), .Y(n29328) );
  INVX1 U17279 ( .A(n33556), .Y(n29335) );
  INVX1 U17280 ( .A(n32190), .Y(n33556) );
  INVX1 U17281 ( .A(n29690), .Y(n34573) );
  INVX1 U17282 ( .A(n32462), .Y(n29329) );
  INVX1 U17283 ( .A(n29668), .Y(n34583) );
  INVX1 U17284 ( .A(n30623), .Y(n30628) );
  INVX1 U17285 ( .A(n30037), .Y(n30622) );
  INVX1 U17286 ( .A(n29339), .Y(n29336) );
  INVX1 U17287 ( .A(n29339), .Y(n29337) );
  INVX1 U17288 ( .A(n29342), .Y(n29340) );
  INVX1 U17289 ( .A(n30471), .Y(n29218) );
  INVX1 U17290 ( .A(n29215), .Y(n29213) );
  INVX1 U17291 ( .A(n30050), .Y(n29215) );
  INVX1 U17292 ( .A(n30050), .Y(n29216) );
  INVX1 U17293 ( .A(n29342), .Y(n29341) );
  INVX1 U17294 ( .A(n29339), .Y(n29338) );
  INVX1 U17295 ( .A(n33059), .Y(n33060) );
  INVX1 U17296 ( .A(n34233), .Y(n34232) );
  INVX1 U17297 ( .A(n34374), .Y(n34375) );
  INVX1 U17298 ( .A(RO[179]), .Y(n32970) );
  INVX1 U17299 ( .A(n3135), .Y(n32811) );
  INVX1 U17300 ( .A(n3130), .Y(n32619) );
  INVX1 U17301 ( .A(n3134), .Y(n32714) );
  INVX1 U17302 ( .A(n3131), .Y(n33010) );
  INVX1 U17303 ( .A(RO[175]), .Y(n32809) );
  INVX1 U17304 ( .A(n3147), .Y(n32883) );
  INVX1 U17305 ( .A(n3171), .Y(n32872) );
  INVX1 U17306 ( .A(n3226), .Y(n32636) );
  INVX1 U17307 ( .A(n3120), .Y(n32677) );
  INVX1 U17308 ( .A(n3121), .Y(n32772) );
  INVX1 U17309 ( .A(oc[0]), .Y(n29755) );
  INVX1 U17310 ( .A(n3154), .Y(n32694) );
  INVX1 U17311 ( .A(n3155), .Y(n32791) );
  INVX1 U17312 ( .A(n3270), .Y(n32584) );
  INVX1 U17313 ( .A(n3271), .Y(n32966) );
  INVX1 U17314 ( .A(n3250), .Y(n32675) );
  INVX1 U17315 ( .A(n3251), .Y(n32769) );
  INVX1 U17316 ( .A(n3184), .Y(n32685) );
  INVX1 U17317 ( .A(n3185), .Y(n32782) );
  INVX1 U17318 ( .A(n12034), .Y(n33389) );
  INVX1 U17319 ( .A(n12066), .Y(n33229) );
  INVX1 U17320 ( .A(n12064), .Y(n33237) );
  INVX1 U17321 ( .A(n12048), .Y(n33321) );
  INVX1 U17322 ( .A(n12046), .Y(n33329) );
  INVX1 U17323 ( .A(n12042), .Y(n33352) );
  INVX1 U17324 ( .A(n12040), .Y(n33359) );
  INVX1 U17325 ( .A(n12028), .Y(n33420) );
  INVX1 U17326 ( .A(n12072), .Y(n33199) );
  INVX1 U17327 ( .A(n12070), .Y(n33206) );
  INVX1 U17328 ( .A(n12076), .Y(n34286) );
  INVX1 U17329 ( .A(n3173), .Y(n32854) );
  INVX1 U17330 ( .A(n3174), .Y(n32667) );
  INVX1 U17331 ( .A(n3175), .Y(n32760) );
  INVX1 U17332 ( .A(n3182), .Y(n32627) );
  INVX1 U17333 ( .A(n3183), .Y(n33018) );
  INVX1 U17334 ( .A(n3202), .Y(n32535) );
  INVX1 U17335 ( .A(n3275), .Y(n32901) );
  INVX1 U17336 ( .A(RO[174]), .Y(n32712) );
  INVX1 U17337 ( .A(n3274), .Y(n32523) );
  INVX1 U17338 ( .A(n3196), .Y(n32648) );
  INVX1 U17339 ( .A(n3198), .Y(n32556) );
  INVX1 U17340 ( .A(n3125), .Y(n32853) );
  INVX1 U17341 ( .A(n3122), .Y(n32573) );
  INVX1 U17342 ( .A(n3126), .Y(n32665) );
  INVX1 U17343 ( .A(n3123), .Y(n32949) );
  INVX1 U17344 ( .A(n3127), .Y(n32758) );
  INVX1 U17345 ( .A(n3160), .Y(n32646) );
  INVX1 U17346 ( .A(n3142), .Y(n32468) );
  INVX1 U17347 ( .A(oc[17]), .Y(n29614) );
  INVX1 U17348 ( .A(oc[23]), .Y(n29612) );
  INVX1 U17349 ( .A(oc[24]), .Y(n29604) );
  INVX1 U17350 ( .A(oc[6]), .Y(n29713) );
  INVX1 U17351 ( .A(RO[178]), .Y(n32587) );
  INVX1 U17352 ( .A(oc[4]), .Y(n29706) );
  XNOR2X1 U17353 ( .A(n23106), .B(n2256), .Y(n27317) );
  XNOR2X1 U17354 ( .A(n27084), .B(n2254), .Y(n27319) );
  XNOR2X1 U17355 ( .A(n25331), .B(n2256), .Y(n27320) );
  XNOR2X1 U17356 ( .A(n25407), .B(n2256), .Y(n27321) );
  INVX1 U17357 ( .A(direct[0]), .Y(n29558) );
  INVX1 U17358 ( .A(n34361), .Y(n34354) );
  AND2X1 U17359 ( .A(invdirect_s2[0]), .B(n33993), .Y(n30663) );
  INVX1 U17360 ( .A(direct[1]), .Y(n29559) );
  INVX1 U17361 ( .A(n3273), .Y(n34225) );
  INVX1 U17362 ( .A(n3272), .Y(n33185) );
  INVX1 U17363 ( .A(n3230), .Y(n33403) );
  INVX1 U17364 ( .A(n3266), .Y(n33220) );
  INVX1 U17365 ( .A(n3267), .Y(n33211) );
  INVX1 U17366 ( .A(n3231), .Y(n33394) );
  INVX1 U17367 ( .A(n3164), .Y(n32740) );
  INVX1 U17368 ( .A(n3114), .Y(n32659) );
  INVX1 U17369 ( .A(n3204), .Y(n32722) );
  INVX1 U17370 ( .A(n3132), .Y(n32602) );
  INVX1 U17371 ( .A(n3162), .Y(n32593) );
  INVX1 U17372 ( .A(n3113), .Y(n32848) );
  INVX1 U17373 ( .A(n3239), .Y(n32912) );
  INVX1 U17374 ( .A(n3112), .Y(n32696) );
  INVX1 U17375 ( .A(n3229), .Y(n32963) );
  INVX1 U17376 ( .A(n3165), .Y(n32952) );
  INVX1 U17377 ( .A(n3115), .Y(n32897) );
  INVX1 U17378 ( .A(n3237), .Y(n33364) );
  INVX1 U17379 ( .A(n3236), .Y(n33373) );
  INVX1 U17380 ( .A(n3228), .Y(n32582) );
  INVX1 U17381 ( .A(n3238), .Y(n32687) );
  INVX1 U17382 ( .A(n3110), .Y(n32567) );
  INVX1 U17383 ( .A(n3111), .Y(n32942) );
  INVX1 U17384 ( .A(address[3]), .Y(n29469) );
  INVX1 U17385 ( .A(n3263), .Y(n33031) );
  INVX1 U17386 ( .A(n3227), .Y(n33029) );
  INVX1 U17387 ( .A(n3170), .Y(n32496) );
  INVX1 U17388 ( .A(n3200), .Y(n32742) );
  INVX1 U17389 ( .A(n3108), .Y(n32604) );
  INVX1 U17390 ( .A(n3144), .Y(n32661) );
  INVX1 U17391 ( .A(n3124), .Y(n32472) );
  INVX1 U17392 ( .A(n3172), .Y(n32474) );
  INVX1 U17393 ( .A(n3141), .Y(n32944) );
  INVX1 U17394 ( .A(n3265), .Y(n32922) );
  INVX1 U17395 ( .A(n3262), .Y(n32638) );
  INVX1 U17396 ( .A(n3201), .Y(n32837) );
  INVX1 U17397 ( .A(n25751), .Y(n32990) );
  INVX1 U17398 ( .A(n3140), .Y(n32569) );
  INVX1 U17399 ( .A(n3264), .Y(n32546) );
  INVX1 U17400 ( .A(n3116), .Y(n32708) );
  INVX1 U17401 ( .A(n3240), .Y(n32724) );
  INVX1 U17402 ( .A(n3241), .Y(n32820) );
  INVX1 U17403 ( .A(n3146), .Y(n32506) );
  INVX1 U17404 ( .A(n3117), .Y(n32805) );
  INVX1 U17405 ( .A(n3248), .Y(n33312) );
  INVX1 U17406 ( .A(n3205), .Y(n32980) );
  INVX1 U17407 ( .A(n3133), .Y(n32987) );
  INVX1 U17408 ( .A(n3163), .Y(n32977) );
  INVX1 U17409 ( .A(n3249), .Y(n33303) );
  INVX1 U17410 ( .A(n3207), .Y(n32874) );
  INVX1 U17411 ( .A(n3206), .Y(n32498) );
  INVX1 U17412 ( .A(n3203), .Y(n32909) );
  INVX1 U17413 ( .A(n3197), .Y(n33040) );
  INVX1 U17414 ( .A(n3145), .Y(n32754) );
  INVX1 U17415 ( .A(n3199), .Y(n32931) );
  INVX1 U17416 ( .A(n3161), .Y(n33038) );
  INVX1 U17417 ( .A(direct[2]), .Y(n29560) );
  INVX1 U17418 ( .A(n3259), .Y(n32803) );
  AND2X2 U17419 ( .A(oc[0]), .B(oc[1]), .Y(n27322) );
  OR2X1 U17420 ( .A(n32571), .B(n32570), .Y(n32577) );
  INVX1 U17421 ( .A(n3257), .Y(n32894) );
  INVX1 U17422 ( .A(n3258), .Y(n32706) );
  OR2X1 U17423 ( .A(n32521), .B(n32520), .Y(n32527) );
  INVX1 U17424 ( .A(n3256), .Y(n32517) );
  INVX1 U17425 ( .A(n3143), .Y(n32850) );
  OR2X1 U17426 ( .A(n32663), .B(n32662), .Y(n32670) );
  INVX1 U17427 ( .A(n30054), .Y(n29192) );
  INVX1 U17428 ( .A(n21151), .Y(n29601) );
  INVX1 U17429 ( .A(wT), .Y(n29526) );
  OR2X1 U17430 ( .A(nc[26]), .B(nc[27]), .Y(n29536) );
  INVX1 U17431 ( .A(nc[6]), .Y(n29542) );
  INVX1 U17432 ( .A(n2254), .Y(n29188) );
  INVX1 U17433 ( .A(S[0]), .Y(n32184) );
  INVX1 U17434 ( .A(nc[16]), .Y(n29531) );
  INVX1 U17435 ( .A(nc[31]), .Y(n29555) );
  INVX1 U17436 ( .A(locTrig[0]), .Y(n30054) );
  INVX1 U17437 ( .A(n8193), .Y(n34134) );
  INVX1 U17438 ( .A(n8194), .Y(n34135) );
  INVX1 U17439 ( .A(n8195), .Y(n34136) );
  INVX1 U17440 ( .A(n8196), .Y(n34137) );
  INVX1 U17441 ( .A(n8197), .Y(n34138) );
  INVX1 U17442 ( .A(n8198), .Y(n34139) );
  INVX1 U17443 ( .A(n8199), .Y(n34140) );
  INVX1 U17444 ( .A(n8200), .Y(n34141) );
  INVX1 U17445 ( .A(n8201), .Y(n34142) );
  INVX1 U17446 ( .A(n8202), .Y(n34143) );
  INVX1 U17447 ( .A(n8203), .Y(n34144) );
  INVX1 U17448 ( .A(n8204), .Y(n34145) );
  INVX1 U17449 ( .A(n8205), .Y(n34146) );
  INVX1 U17450 ( .A(n8206), .Y(n34147) );
  INVX1 U17451 ( .A(n8207), .Y(n34148) );
  INVX1 U17452 ( .A(n8208), .Y(n34149) );
  INVX1 U17453 ( .A(n8209), .Y(n34150) );
  INVX1 U17454 ( .A(n8210), .Y(n34151) );
  INVX1 U17455 ( .A(n8211), .Y(n34152) );
  INVX1 U17456 ( .A(n8212), .Y(n34153) );
  INVX1 U17457 ( .A(n8213), .Y(n34154) );
  INVX1 U17458 ( .A(n8214), .Y(n34155) );
  INVX1 U17459 ( .A(n8215), .Y(n34156) );
  INVX1 U17460 ( .A(n8216), .Y(n34157) );
  INVX1 U17461 ( .A(n8217), .Y(n34158) );
  INVX1 U17462 ( .A(n8218), .Y(n34159) );
  INVX1 U17463 ( .A(n8154), .Y(n34095) );
  INVX1 U17464 ( .A(n8155), .Y(n34096) );
  INVX1 U17465 ( .A(n8156), .Y(n34097) );
  INVX1 U17466 ( .A(n8157), .Y(n34098) );
  INVX1 U17467 ( .A(n8158), .Y(n34099) );
  INVX1 U17468 ( .A(n8159), .Y(n34100) );
  INVX1 U17469 ( .A(n8160), .Y(n34101) );
  INVX1 U17470 ( .A(n8161), .Y(n34102) );
  INVX1 U17471 ( .A(n8162), .Y(n34103) );
  INVX1 U17472 ( .A(n8163), .Y(n34104) );
  INVX1 U17473 ( .A(n8164), .Y(n34105) );
  INVX1 U17474 ( .A(n8165), .Y(n34106) );
  INVX1 U17475 ( .A(n8166), .Y(n34107) );
  INVX1 U17476 ( .A(n8167), .Y(n34108) );
  INVX1 U17477 ( .A(n8168), .Y(n34109) );
  INVX1 U17478 ( .A(n8169), .Y(n34110) );
  INVX1 U17479 ( .A(n8170), .Y(n34111) );
  INVX1 U17480 ( .A(n8171), .Y(n34112) );
  INVX1 U17481 ( .A(n8172), .Y(n34113) );
  INVX1 U17482 ( .A(n8173), .Y(n34114) );
  INVX1 U17483 ( .A(n8174), .Y(n34115) );
  INVX1 U17484 ( .A(n8175), .Y(n34116) );
  INVX1 U17485 ( .A(n8176), .Y(n34117) );
  INVX1 U17486 ( .A(n8177), .Y(n34118) );
  INVX1 U17487 ( .A(n8178), .Y(n34119) );
  INVX1 U17488 ( .A(n8179), .Y(n34120) );
  INVX1 U17489 ( .A(n8180), .Y(n34121) );
  INVX1 U17490 ( .A(n8181), .Y(n34122) );
  INVX1 U17491 ( .A(n8182), .Y(n34123) );
  INVX1 U17492 ( .A(n8183), .Y(n34124) );
  INVX1 U17493 ( .A(n8184), .Y(n34125) );
  INVX1 U17494 ( .A(n8185), .Y(n34126) );
  INVX1 U17495 ( .A(n8186), .Y(n34127) );
  INVX1 U17496 ( .A(n8187), .Y(n34128) );
  INVX1 U17497 ( .A(n8188), .Y(n34129) );
  INVX1 U17498 ( .A(n8189), .Y(n34130) );
  INVX1 U17499 ( .A(n8190), .Y(n34131) );
  INVX1 U17500 ( .A(n8191), .Y(n34132) );
  INVX1 U17501 ( .A(n8192), .Y(n34133) );
  INVX1 U17502 ( .A(n8219), .Y(n34160) );
  INVX1 U17503 ( .A(n8220), .Y(n34161) );
  INVX1 U17504 ( .A(n8221), .Y(n34162) );
  INVX1 U17505 ( .A(n8222), .Y(n34163) );
  INVX1 U17506 ( .A(n8223), .Y(n34164) );
  INVX1 U17507 ( .A(n8224), .Y(n34165) );
  INVX1 U17508 ( .A(n8225), .Y(n34166) );
  INVX1 U17509 ( .A(n8226), .Y(n34167) );
  INVX1 U17510 ( .A(n8227), .Y(n34168) );
  INVX1 U17511 ( .A(n8228), .Y(n34169) );
  INVX1 U17512 ( .A(n8229), .Y(n34229) );
  INVX1 U17513 ( .A(n8076), .Y(n34017) );
  INVX1 U17514 ( .A(n8077), .Y(n34018) );
  INVX1 U17515 ( .A(n8078), .Y(n34019) );
  INVX1 U17516 ( .A(n8079), .Y(n34020) );
  INVX1 U17517 ( .A(n8080), .Y(n34021) );
  INVX1 U17518 ( .A(n8081), .Y(n34022) );
  INVX1 U17519 ( .A(n8082), .Y(n34023) );
  INVX1 U17520 ( .A(n8083), .Y(n34024) );
  INVX1 U17521 ( .A(n8084), .Y(n34025) );
  INVX1 U17522 ( .A(n8085), .Y(n34026) );
  INVX1 U17523 ( .A(n8086), .Y(n34027) );
  INVX1 U17524 ( .A(n8087), .Y(n34028) );
  INVX1 U17525 ( .A(n8088), .Y(n34029) );
  INVX1 U17526 ( .A(n8089), .Y(n34030) );
  INVX1 U17527 ( .A(n8090), .Y(n34031) );
  INVX1 U17528 ( .A(n8091), .Y(n34032) );
  INVX1 U17529 ( .A(n8092), .Y(n34033) );
  INVX1 U17530 ( .A(n8093), .Y(n34034) );
  INVX1 U17531 ( .A(n8094), .Y(n34035) );
  INVX1 U17532 ( .A(n8095), .Y(n34036) );
  INVX1 U17533 ( .A(n8096), .Y(n34037) );
  INVX1 U17534 ( .A(n8097), .Y(n34038) );
  INVX1 U17535 ( .A(n8098), .Y(n34039) );
  INVX1 U17536 ( .A(n8099), .Y(n34040) );
  INVX1 U17537 ( .A(n8100), .Y(n34041) );
  INVX1 U17538 ( .A(n8101), .Y(n34042) );
  INVX1 U17539 ( .A(n8102), .Y(n34043) );
  INVX1 U17540 ( .A(n8103), .Y(n34044) );
  INVX1 U17541 ( .A(n8104), .Y(n34045) );
  INVX1 U17542 ( .A(n8105), .Y(n34046) );
  INVX1 U17543 ( .A(n8106), .Y(n34047) );
  INVX1 U17544 ( .A(n8107), .Y(n34048) );
  INVX1 U17545 ( .A(n8108), .Y(n34049) );
  INVX1 U17546 ( .A(n8109), .Y(n34050) );
  INVX1 U17547 ( .A(n8110), .Y(n34051) );
  INVX1 U17548 ( .A(n8111), .Y(n34052) );
  INVX1 U17549 ( .A(n8112), .Y(n34053) );
  INVX1 U17550 ( .A(n8113), .Y(n34054) );
  INVX1 U17551 ( .A(n8114), .Y(n34055) );
  INVX1 U17552 ( .A(n8115), .Y(n34056) );
  INVX1 U17553 ( .A(n8116), .Y(n34057) );
  INVX1 U17554 ( .A(n8117), .Y(n34058) );
  INVX1 U17555 ( .A(n8118), .Y(n34059) );
  INVX1 U17556 ( .A(n8119), .Y(n34060) );
  INVX1 U17557 ( .A(n8120), .Y(n34061) );
  INVX1 U17558 ( .A(n8121), .Y(n34062) );
  INVX1 U17559 ( .A(n8122), .Y(n34063) );
  INVX1 U17560 ( .A(n8123), .Y(n34064) );
  INVX1 U17561 ( .A(n8124), .Y(n34065) );
  INVX1 U17562 ( .A(n8125), .Y(n34066) );
  INVX1 U17563 ( .A(n8126), .Y(n34067) );
  INVX1 U17564 ( .A(n8127), .Y(n34068) );
  INVX1 U17565 ( .A(n8128), .Y(n34069) );
  INVX1 U17566 ( .A(n8129), .Y(n34070) );
  INVX1 U17567 ( .A(n8130), .Y(n34071) );
  INVX1 U17568 ( .A(n8131), .Y(n34072) );
  INVX1 U17569 ( .A(n8132), .Y(n34073) );
  INVX1 U17570 ( .A(n8133), .Y(n34074) );
  INVX1 U17571 ( .A(n8134), .Y(n34075) );
  INVX1 U17572 ( .A(n8135), .Y(n34076) );
  INVX1 U17573 ( .A(n8136), .Y(n34077) );
  INVX1 U17574 ( .A(n8137), .Y(n34078) );
  INVX1 U17575 ( .A(n8138), .Y(n34079) );
  INVX1 U17576 ( .A(n8139), .Y(n34080) );
  INVX1 U17577 ( .A(n8140), .Y(n34081) );
  INVX1 U17578 ( .A(n8141), .Y(n34082) );
  INVX1 U17579 ( .A(n8142), .Y(n34083) );
  INVX1 U17580 ( .A(n8143), .Y(n34084) );
  INVX1 U17581 ( .A(n8144), .Y(n34085) );
  INVX1 U17582 ( .A(n8145), .Y(n34086) );
  INVX1 U17583 ( .A(n8146), .Y(n34087) );
  INVX1 U17584 ( .A(n8147), .Y(n34088) );
  INVX1 U17585 ( .A(n8148), .Y(n34089) );
  INVX1 U17586 ( .A(n8149), .Y(n34090) );
  INVX1 U17587 ( .A(n8150), .Y(n34091) );
  INVX1 U17588 ( .A(n8151), .Y(n34092) );
  INVX1 U17589 ( .A(n8152), .Y(n34093) );
  INVX1 U17590 ( .A(n8153), .Y(n34094) );
  INVX1 U17591 ( .A(n8056), .Y(n33997) );
  INVX1 U17592 ( .A(n8057), .Y(n33998) );
  INVX1 U17593 ( .A(n8058), .Y(n33999) );
  INVX1 U17594 ( .A(n8059), .Y(n34000) );
  INVX1 U17595 ( .A(n8060), .Y(n34001) );
  INVX1 U17596 ( .A(n8061), .Y(n34002) );
  INVX1 U17597 ( .A(n8062), .Y(n34003) );
  INVX1 U17598 ( .A(n8063), .Y(n34004) );
  INVX1 U17599 ( .A(n8064), .Y(n34005) );
  INVX1 U17600 ( .A(n8065), .Y(n34006) );
  INVX1 U17601 ( .A(n8066), .Y(n34007) );
  INVX1 U17602 ( .A(n8067), .Y(n34008) );
  INVX1 U17603 ( .A(n8068), .Y(n34009) );
  INVX1 U17604 ( .A(n8069), .Y(n34010) );
  INVX1 U17605 ( .A(n8070), .Y(n34011) );
  INVX1 U17606 ( .A(n8071), .Y(n34012) );
  INVX1 U17607 ( .A(n8072), .Y(n34013) );
  INVX1 U17608 ( .A(n8073), .Y(n34014) );
  INVX1 U17609 ( .A(n8074), .Y(n34015) );
  INVX1 U17610 ( .A(n8075), .Y(n34016) );
  INVX1 U17611 ( .A(nc[2]), .Y(n29550) );
  INVX1 U17612 ( .A(nc[20]), .Y(n29528) );
  INVX1 U17613 ( .A(nc[21]), .Y(n29530) );
  INVX1 U17614 ( .A(nc[17]), .Y(n29533) );
  INVX1 U17615 ( .A(n30074), .Y(n30643) );
  INVX1 U17616 ( .A(n34283), .Y(n29404) );
  INVX1 U17617 ( .A(n34341), .Y(n29413) );
  INVX1 U17618 ( .A(n34343), .Y(n29421) );
  INVX1 U17619 ( .A(n3255), .Y(n33272) );
  INVX1 U17620 ( .A(n3254), .Y(n33281) );
  INVX1 U17621 ( .A(n3225), .Y(n33425) );
  INVX1 U17622 ( .A(n3242), .Y(n33343) );
  INVX1 U17623 ( .A(n3243), .Y(n33334) );
  INVX1 U17624 ( .A(Setup[0]), .Y(n29703) );
  INVX1 U17625 ( .A(n3260), .Y(n33251) );
  INVX1 U17626 ( .A(n3261), .Y(n33242) );
  INVX1 U17627 ( .A(states[1]), .Y(n29603) );
  INVX1 U17628 ( .A(states[0]), .Y(n29527) );
  INVX1 U17629 ( .A(n34282), .Y(n29395) );
  INVX1 U17630 ( .A(T[1]), .Y(n34372) );
  AND2X1 U17631 ( .A(n15177), .B(data_in[0]), .Y(n27323) );
  AND2X1 U17632 ( .A(data_in[4]), .B(n15174), .Y(n27324) );
  INVX1 U17633 ( .A(n30235), .Y(n30272) );
  INVX1 U17634 ( .A(n30372), .Y(n30409) );
  INVX1 U17635 ( .A(n30185), .Y(n30225) );
  INVX1 U17636 ( .A(n30280), .Y(n30319) );
  INVX1 U17637 ( .A(n30143), .Y(n30179) );
  INVX1 U17638 ( .A(n30101), .Y(n30440) );
  INVX1 U17639 ( .A(n30118), .Y(n30457) );
  INVX1 U17640 ( .A(n30085), .Y(n30426) );
  INVX1 U17641 ( .A(n30092), .Y(n30432) );
  INVX1 U17642 ( .A(n30109), .Y(n30449) );
  INVX1 U17643 ( .A(T[0]), .Y(n34379) );
  AND2X1 U17644 ( .A(data_in[2]), .B(data_in[1]), .Y(n15177) );
  INVX1 U17645 ( .A(data_in[4]), .Y(n30327) );
  INVX1 U17646 ( .A(data_in[0]), .Y(n30126) );
  INVX1 U17647 ( .A(data_in[5]), .Y(n30234) );
  INVX1 U17648 ( .A(data_in[2]), .Y(n30100) );
  INVX1 U17649 ( .A(data_in[1]), .Y(n30117) );
  INVX1 U17650 ( .A(data_in[3]), .Y(n30371) );
  INVX1 U17651 ( .A(T[4]), .Y(n34356) );
  INVX1 U17652 ( .A(T[5]), .Y(n34351) );
  INVX1 U17653 ( .A(T[3]), .Y(n34360) );
  INVX1 U17654 ( .A(T[2]), .Y(n34385) );
  INVX1 U17655 ( .A(S[5]), .Y(n32159) );
  INVX1 U17656 ( .A(S[4]), .Y(n32164) );
  INVX1 U17657 ( .A(S[3]), .Y(n32169) );
  INVX1 U17658 ( .A(S[2]), .Y(n32174) );
  INVX1 U17659 ( .A(S[1]), .Y(n32179) );
  INVX1 U17660 ( .A(n29681), .Y(n29682) );
  INVX1 U17661 ( .A(n29648), .Y(n29640) );
  INVX1 U17662 ( .A(n20812), .Y(n34615) );
  INVX1 U17663 ( .A(n29677), .Y(n29675) );
  INVX1 U17664 ( .A(n29671), .Y(n29669) );
  INVX1 U17665 ( .A(n29651), .Y(n29650) );
  INVX1 U17666 ( .A(n29659), .Y(n29658) );
  XNOR2X1 U17667 ( .A(n23611), .B(T[1]), .Y(n27325) );
  INVX1 U17668 ( .A(n14870), .Y(n34607) );
  INVX1 U17669 ( .A(n14673), .Y(n34610) );
  INVX1 U17670 ( .A(n14575), .Y(n34600) );
  INVX1 U17671 ( .A(n29688), .Y(n29689) );
  INVX1 U17672 ( .A(n29666), .Y(n29667) );
  INVX1 U17673 ( .A(n14477), .Y(n34604) );
  INVX1 U17674 ( .A(address[5]), .Y(n34616) );
  INVX1 U17675 ( .A(n16149), .Y(n34556) );
  INVX1 U17676 ( .A(n32193), .Y(n32462) );
  XNOR2X1 U17677 ( .A(n29666), .B(T[1]), .Y(n27326) );
  XNOR2X1 U17678 ( .A(n29688), .B(T[1]), .Y(n27327) );
  OR2X1 U17679 ( .A(n15182), .B(n15183), .Y(n30070) );
  INVX1 U17680 ( .A(Setup[1]), .Y(n34505) );
  INVX1 U17681 ( .A(n33557), .Y(n29339) );
  INVX1 U17682 ( .A(n30488), .Y(n33557) );
  OR2X1 U17683 ( .A(n2266), .B(n2265), .Y(n15178) );
  INVX1 U17684 ( .A(wS), .Y(n34614) );
  INVX1 U17685 ( .A(n33559), .Y(n29342) );
  INVX1 U17686 ( .A(n30490), .Y(n33559) );
  INVX1 U17687 ( .A(addrLock), .Y(n30067) );
  INVX1 U17688 ( .A(n14354), .Y(n13743) );
  INVX1 U17689 ( .A(n33174), .Y(n22636) );
  INVX1 U17690 ( .A(n29895), .Y(n15544) );
  INVX1 U17691 ( .A(n29889), .Y(n15552) );
  OR2X1 U17692 ( .A(n15580), .B(n14218), .Y(n22372) );
  INVX1 U17693 ( .A(n30550), .Y(n30554) );
  INVX1 U17694 ( .A(n15873), .Y(n29740) );
  INVX1 U17695 ( .A(n22323), .Y(n13994) );
  MUX2X1 U17696 ( .B(n27329), .A(n27330), .S(n27701), .Y(n27328) );
  MUX2X1 U17697 ( .B(n27332), .A(n27333), .S(n27701), .Y(n27331) );
  MUX2X1 U17698 ( .B(n27335), .A(n27336), .S(n27701), .Y(n27334) );
  MUX2X1 U17699 ( .B(n27338), .A(n27339), .S(n27701), .Y(n27337) );
  MUX2X1 U17700 ( .B(n27341), .A(n27342), .S(n27704), .Y(n27340) );
  MUX2X1 U17701 ( .B(n27344), .A(n27345), .S(n27701), .Y(n27343) );
  MUX2X1 U17702 ( .B(n27347), .A(n27348), .S(n27701), .Y(n27346) );
  MUX2X1 U17703 ( .B(n27350), .A(n27351), .S(n27701), .Y(n27349) );
  MUX2X1 U17704 ( .B(n27353), .A(n27354), .S(n27701), .Y(n27352) );
  MUX2X1 U17705 ( .B(n27356), .A(n27357), .S(n27704), .Y(n27355) );
  MUX2X1 U17706 ( .B(n27359), .A(n27360), .S(n27701), .Y(n27358) );
  MUX2X1 U17707 ( .B(n27362), .A(n27363), .S(n27701), .Y(n27361) );
  MUX2X1 U17708 ( .B(n27365), .A(n27366), .S(n27701), .Y(n27364) );
  MUX2X1 U17709 ( .B(n27368), .A(n27369), .S(n27701), .Y(n27367) );
  MUX2X1 U17710 ( .B(n27371), .A(n27372), .S(n27704), .Y(n27370) );
  MUX2X1 U17711 ( .B(n27374), .A(n27375), .S(n27701), .Y(n27373) );
  MUX2X1 U17712 ( .B(n27377), .A(n27378), .S(n27700), .Y(n27376) );
  MUX2X1 U17713 ( .B(n27380), .A(n27381), .S(n27701), .Y(n27379) );
  MUX2X1 U17714 ( .B(n27383), .A(n27384), .S(n27700), .Y(n27382) );
  MUX2X1 U17715 ( .B(n27386), .A(n27387), .S(n27704), .Y(n27385) );
  MUX2X1 U17716 ( .B(n27388), .A(n27389), .S(n20975), .Y(n2266) );
  MUX2X1 U17717 ( .B(n27391), .A(n27392), .S(n27700), .Y(n27390) );
  MUX2X1 U17718 ( .B(n27394), .A(n27395), .S(n27700), .Y(n27393) );
  MUX2X1 U17719 ( .B(n27397), .A(n27398), .S(n27701), .Y(n27396) );
  MUX2X1 U17720 ( .B(n27400), .A(n27401), .S(n27700), .Y(n27399) );
  MUX2X1 U17721 ( .B(n27403), .A(n27404), .S(n27704), .Y(n27402) );
  MUX2X1 U17722 ( .B(n27406), .A(n27407), .S(n27700), .Y(n27405) );
  MUX2X1 U17723 ( .B(n27409), .A(n27410), .S(n27700), .Y(n27408) );
  MUX2X1 U17724 ( .B(n27412), .A(n27413), .S(n27701), .Y(n27411) );
  MUX2X1 U17725 ( .B(n27415), .A(n27416), .S(n27701), .Y(n27414) );
  MUX2X1 U17726 ( .B(n27418), .A(n27419), .S(n27704), .Y(n27417) );
  MUX2X1 U17727 ( .B(n27421), .A(n27422), .S(n27700), .Y(n27420) );
  MUX2X1 U17728 ( .B(n27424), .A(n27425), .S(n27700), .Y(n27423) );
  MUX2X1 U17729 ( .B(n27427), .A(n27428), .S(n27700), .Y(n27426) );
  MUX2X1 U17730 ( .B(n27430), .A(n27431), .S(n27700), .Y(n27429) );
  MUX2X1 U17731 ( .B(n27433), .A(n27434), .S(n27704), .Y(n27432) );
  MUX2X1 U17732 ( .B(n27436), .A(n27437), .S(n27700), .Y(n27435) );
  MUX2X1 U17733 ( .B(n27439), .A(n27440), .S(n27700), .Y(n27438) );
  MUX2X1 U17734 ( .B(n27442), .A(n27443), .S(n27700), .Y(n27441) );
  MUX2X1 U17735 ( .B(n27445), .A(n27446), .S(n27700), .Y(n27444) );
  MUX2X1 U17736 ( .B(n27448), .A(n27449), .S(n27704), .Y(n27447) );
  MUX2X1 U17737 ( .B(n27450), .A(n27451), .S(n20975), .Y(n2265) );
  MUX2X1 U17738 ( .B(n27453), .A(n27454), .S(n27700), .Y(n27452) );
  MUX2X1 U17739 ( .B(n27456), .A(n27457), .S(n27700), .Y(n27455) );
  MUX2X1 U17740 ( .B(n27459), .A(n27460), .S(n27700), .Y(n27458) );
  MUX2X1 U17741 ( .B(n27462), .A(n27463), .S(n27700), .Y(n27461) );
  MUX2X1 U17742 ( .B(n27465), .A(n27466), .S(n27704), .Y(n27464) );
  MUX2X1 U17743 ( .B(n27468), .A(n27469), .S(n27701), .Y(n27467) );
  MUX2X1 U17744 ( .B(n27471), .A(n27472), .S(n27700), .Y(n27470) );
  MUX2X1 U17745 ( .B(n27474), .A(n27475), .S(n27701), .Y(n27473) );
  MUX2X1 U17746 ( .B(n27477), .A(n27478), .S(n27700), .Y(n27476) );
  MUX2X1 U17747 ( .B(n27480), .A(n27481), .S(n27704), .Y(n27479) );
  MUX2X1 U17748 ( .B(n27483), .A(n27484), .S(n27701), .Y(n27482) );
  MUX2X1 U17749 ( .B(n27486), .A(n27487), .S(n27700), .Y(n27485) );
  MUX2X1 U17750 ( .B(n27489), .A(n27490), .S(n27701), .Y(n27488) );
  MUX2X1 U17751 ( .B(n27492), .A(n27493), .S(n27700), .Y(n27491) );
  MUX2X1 U17752 ( .B(n27495), .A(n27496), .S(n27704), .Y(n27494) );
  MUX2X1 U17753 ( .B(n27498), .A(n27499), .S(n27701), .Y(n27497) );
  MUX2X1 U17754 ( .B(n27501), .A(n27502), .S(n27700), .Y(n27500) );
  MUX2X1 U17755 ( .B(n27504), .A(n27505), .S(n27701), .Y(n27503) );
  MUX2X1 U17756 ( .B(n27507), .A(n27508), .S(n27700), .Y(n27506) );
  MUX2X1 U17757 ( .B(n27510), .A(n27511), .S(n27704), .Y(n27509) );
  MUX2X1 U17758 ( .B(n27512), .A(n27513), .S(n20975), .Y(n2264) );
  MUX2X1 U17759 ( .B(n27515), .A(n27516), .S(n27701), .Y(n27514) );
  MUX2X1 U17760 ( .B(n27518), .A(n27519), .S(n27701), .Y(n27517) );
  MUX2X1 U17761 ( .B(n27521), .A(n27522), .S(n27700), .Y(n27520) );
  MUX2X1 U17762 ( .B(n27524), .A(n27525), .S(n27701), .Y(n27523) );
  MUX2X1 U17763 ( .B(n27527), .A(n27528), .S(n27704), .Y(n27526) );
  MUX2X1 U17764 ( .B(n27530), .A(n27531), .S(n27700), .Y(n27529) );
  MUX2X1 U17765 ( .B(n27533), .A(n27534), .S(n27700), .Y(n27532) );
  MUX2X1 U17766 ( .B(n27536), .A(n27537), .S(n27701), .Y(n27535) );
  MUX2X1 U17767 ( .B(n27539), .A(n27540), .S(n27701), .Y(n27538) );
  MUX2X1 U17768 ( .B(n27542), .A(n27543), .S(n27704), .Y(n27541) );
  MUX2X1 U17769 ( .B(n27545), .A(n27546), .S(n27700), .Y(n27544) );
  MUX2X1 U17770 ( .B(n27548), .A(n27549), .S(n27701), .Y(n27547) );
  MUX2X1 U17771 ( .B(n27551), .A(n27552), .S(n27700), .Y(n27550) );
  MUX2X1 U17772 ( .B(n27554), .A(n27555), .S(n27700), .Y(n27553) );
  MUX2X1 U17773 ( .B(n27557), .A(n27558), .S(n27704), .Y(n27556) );
  MUX2X1 U17774 ( .B(n27560), .A(n27561), .S(n27701), .Y(n27559) );
  MUX2X1 U17775 ( .B(n27563), .A(n27564), .S(n27700), .Y(n27562) );
  MUX2X1 U17776 ( .B(n27566), .A(n27567), .S(n27700), .Y(n27565) );
  MUX2X1 U17777 ( .B(n27569), .A(n27570), .S(n27700), .Y(n27568) );
  MUX2X1 U17778 ( .B(n27572), .A(n27573), .S(n27704), .Y(n27571) );
  MUX2X1 U17779 ( .B(n27574), .A(n27575), .S(n20975), .Y(n2263) );
  MUX2X1 U17780 ( .B(n27577), .A(n27578), .S(n27701), .Y(n27576) );
  MUX2X1 U17781 ( .B(n27580), .A(n27581), .S(n27701), .Y(n27579) );
  MUX2X1 U17782 ( .B(n27583), .A(n27584), .S(n27700), .Y(n27582) );
  MUX2X1 U17783 ( .B(n27586), .A(n27587), .S(n27701), .Y(n27585) );
  MUX2X1 U17784 ( .B(n27589), .A(n27590), .S(n27704), .Y(n27588) );
  MUX2X1 U17785 ( .B(n27592), .A(n27593), .S(n27701), .Y(n27591) );
  MUX2X1 U17786 ( .B(n27595), .A(n27596), .S(n27700), .Y(n27594) );
  MUX2X1 U17787 ( .B(n27598), .A(n27599), .S(n27700), .Y(n27597) );
  MUX2X1 U17788 ( .B(n27601), .A(n27602), .S(n27700), .Y(n27600) );
  MUX2X1 U17789 ( .B(n27604), .A(n27605), .S(n27704), .Y(n27603) );
  MUX2X1 U17790 ( .B(n27607), .A(n27608), .S(n27700), .Y(n27606) );
  MUX2X1 U17791 ( .B(n27610), .A(n27611), .S(n27701), .Y(n27609) );
  MUX2X1 U17792 ( .B(n27613), .A(n27614), .S(n27701), .Y(n27612) );
  MUX2X1 U17793 ( .B(n27616), .A(n27617), .S(n27701), .Y(n27615) );
  MUX2X1 U17794 ( .B(n27619), .A(n27620), .S(n27704), .Y(n27618) );
  MUX2X1 U17795 ( .B(n27622), .A(n27623), .S(n27700), .Y(n27621) );
  MUX2X1 U17796 ( .B(n27625), .A(n27626), .S(n27700), .Y(n27624) );
  MUX2X1 U17797 ( .B(n27628), .A(n27629), .S(n27701), .Y(n27627) );
  MUX2X1 U17798 ( .B(n27631), .A(n27632), .S(n27700), .Y(n27630) );
  MUX2X1 U17799 ( .B(n27634), .A(n27635), .S(n27704), .Y(n27633) );
  MUX2X1 U17800 ( .B(n27636), .A(n27637), .S(n20975), .Y(n2262) );
  MUX2X1 U17801 ( .B(n27639), .A(n27640), .S(n27700), .Y(n27638) );
  MUX2X1 U17802 ( .B(n27642), .A(n27643), .S(n27700), .Y(n27641) );
  MUX2X1 U17803 ( .B(n27645), .A(n27646), .S(n27701), .Y(n27644) );
  MUX2X1 U17804 ( .B(n27648), .A(n27649), .S(n27701), .Y(n27647) );
  MUX2X1 U17805 ( .B(n27651), .A(n27652), .S(n27704), .Y(n27650) );
  MUX2X1 U17806 ( .B(n27654), .A(n27655), .S(n27701), .Y(n27653) );
  MUX2X1 U17807 ( .B(n27657), .A(n27658), .S(n27701), .Y(n27656) );
  MUX2X1 U17808 ( .B(n27660), .A(n27661), .S(n27700), .Y(n27659) );
  MUX2X1 U17809 ( .B(n27663), .A(n27664), .S(n27701), .Y(n27662) );
  MUX2X1 U17810 ( .B(n27666), .A(n27667), .S(n27704), .Y(n27665) );
  MUX2X1 U17811 ( .B(n27669), .A(n27670), .S(n27700), .Y(n27668) );
  MUX2X1 U17812 ( .B(n27672), .A(n27673), .S(n27701), .Y(n27671) );
  MUX2X1 U17813 ( .B(n27675), .A(n27676), .S(n27701), .Y(n27674) );
  MUX2X1 U17814 ( .B(n27678), .A(n27679), .S(n27701), .Y(n27677) );
  MUX2X1 U17815 ( .B(n27681), .A(n27682), .S(n27704), .Y(n27680) );
  MUX2X1 U17816 ( .B(n27684), .A(n27685), .S(n27700), .Y(n27683) );
  MUX2X1 U17817 ( .B(n27687), .A(n27688), .S(n27700), .Y(n27686) );
  MUX2X1 U17818 ( .B(n27690), .A(n27691), .S(n27701), .Y(n27689) );
  MUX2X1 U17819 ( .B(n27693), .A(n27694), .S(n27701), .Y(n27692) );
  MUX2X1 U17820 ( .B(n27696), .A(n27697), .S(n27704), .Y(n27695) );
  MUX2X1 U17821 ( .B(n27698), .A(n27699), .S(n20975), .Y(n2261) );
  MUX2X1 U17822 ( .B(grid[372]), .A(grid[378]), .S(n27714), .Y(n27330) );
  MUX2X1 U17823 ( .B(n21081), .A(grid[366]), .S(n27714), .Y(n27329) );
  MUX2X1 U17824 ( .B(n25626), .A(grid[354]), .S(n27714), .Y(n27333) );
  MUX2X1 U17825 ( .B(grid[336]), .A(grid[342]), .S(n27714), .Y(n27332) );
  MUX2X1 U17826 ( .B(n27331), .A(n27328), .S(n27702), .Y(n27342) );
  MUX2X1 U17827 ( .B(grid[324]), .A(grid[330]), .S(n27714), .Y(n27336) );
  MUX2X1 U17828 ( .B(grid[312]), .A(grid[318]), .S(n27714), .Y(n27335) );
  MUX2X1 U17829 ( .B(n25618), .A(grid[306]), .S(n27714), .Y(n27339) );
  MUX2X1 U17830 ( .B(grid[288]), .A(grid[294]), .S(n27714), .Y(n27338) );
  MUX2X1 U17831 ( .B(n27337), .A(n27334), .S(n27702), .Y(n27341) );
  MUX2X1 U17832 ( .B(n25627), .A(grid[282]), .S(n27714), .Y(n27345) );
  MUX2X1 U17833 ( .B(grid[264]), .A(grid[270]), .S(n27714), .Y(n27344) );
  MUX2X1 U17834 ( .B(n25643), .A(grid[258]), .S(n27714), .Y(n27348) );
  MUX2X1 U17835 ( .B(n25637), .A(grid[246]), .S(n27714), .Y(n27347) );
  MUX2X1 U17836 ( .B(n27346), .A(n27343), .S(n27702), .Y(n27357) );
  MUX2X1 U17837 ( .B(n21088), .A(grid[234]), .S(n27713), .Y(n27351) );
  MUX2X1 U17838 ( .B(grid[216]), .A(grid[222]), .S(n27713), .Y(n27350) );
  MUX2X1 U17839 ( .B(n25635), .A(grid[210]), .S(n27713), .Y(n27354) );
  MUX2X1 U17840 ( .B(n25631), .A(grid[198]), .S(n27713), .Y(n27353) );
  MUX2X1 U17841 ( .B(n27352), .A(n27349), .S(n27702), .Y(n27356) );
  MUX2X1 U17842 ( .B(n27355), .A(n27340), .S(n20812), .Y(n27389) );
  MUX2X1 U17843 ( .B(grid[180]), .A(grid[186]), .S(n27713), .Y(n27360) );
  MUX2X1 U17844 ( .B(grid[168]), .A(grid[174]), .S(n27713), .Y(n27359) );
  MUX2X1 U17845 ( .B(grid[156]), .A(n25625), .S(n27713), .Y(n27363) );
  MUX2X1 U17846 ( .B(n21084), .A(grid[150]), .S(n27713), .Y(n27362) );
  MUX2X1 U17847 ( .B(n27361), .A(n27358), .S(n27702), .Y(n27372) );
  MUX2X1 U17848 ( .B(grid[132]), .A(grid[138]), .S(n27713), .Y(n27366) );
  MUX2X1 U17849 ( .B(grid[120]), .A(grid[126]), .S(n27713), .Y(n27365) );
  MUX2X1 U17850 ( .B(grid[108]), .A(grid[114]), .S(n27713), .Y(n27369) );
  MUX2X1 U17851 ( .B(grid[96]), .A(grid[102]), .S(n27713), .Y(n27368) );
  MUX2X1 U17852 ( .B(n27367), .A(n27364), .S(n27702), .Y(n27371) );
  MUX2X1 U17853 ( .B(grid[84]), .A(n21082), .S(n27712), .Y(n27375) );
  MUX2X1 U17854 ( .B(grid[72]), .A(grid[78]), .S(n27712), .Y(n27374) );
  MUX2X1 U17855 ( .B(n25639), .A(n25478), .S(n27712), .Y(n27378) );
  MUX2X1 U17856 ( .B(n25632), .A(grid[54]), .S(n27712), .Y(n27377) );
  MUX2X1 U17857 ( .B(n27376), .A(n27373), .S(n27702), .Y(n27387) );
  MUX2X1 U17858 ( .B(n21087), .A(grid[42]), .S(n27712), .Y(n27381) );
  MUX2X1 U17859 ( .B(grid[24]), .A(n21083), .S(n27712), .Y(n27380) );
  MUX2X1 U17860 ( .B(n25633), .A(grid[18]), .S(n27712), .Y(n27384) );
  MUX2X1 U17861 ( .B(grid[0]), .A(n21086), .S(n27712), .Y(n27383) );
  MUX2X1 U17862 ( .B(n27382), .A(n27379), .S(n27702), .Y(n27386) );
  MUX2X1 U17863 ( .B(n27385), .A(n27370), .S(n20812), .Y(n27388) );
  MUX2X1 U17864 ( .B(grid[373]), .A(grid[379]), .S(n27712), .Y(n27392) );
  MUX2X1 U17865 ( .B(grid[361]), .A(n21215), .S(n27712), .Y(n27391) );
  MUX2X1 U17866 ( .B(n25488), .A(n25498), .S(n27712), .Y(n27395) );
  MUX2X1 U17867 ( .B(grid[337]), .A(n25492), .S(n27712), .Y(n27394) );
  MUX2X1 U17868 ( .B(n27393), .A(n27390), .S(n27702), .Y(n27404) );
  MUX2X1 U17869 ( .B(grid[325]), .A(n23205), .S(n27711), .Y(n27398) );
  MUX2X1 U17870 ( .B(grid[313]), .A(grid[319]), .S(n27711), .Y(n27397) );
  MUX2X1 U17871 ( .B(n20845), .A(n25493), .S(n27711), .Y(n27401) );
  MUX2X1 U17872 ( .B(grid[289]), .A(grid[295]), .S(n27711), .Y(n27400) );
  MUX2X1 U17873 ( .B(n27399), .A(n27396), .S(n27702), .Y(n27403) );
  MUX2X1 U17874 ( .B(n25583), .A(grid[283]), .S(n27711), .Y(n27407) );
  MUX2X1 U17875 ( .B(n25506), .A(grid[271]), .S(n27711), .Y(n27406) );
  MUX2X1 U17876 ( .B(n25490), .A(grid[259]), .S(n27711), .Y(n27410) );
  MUX2X1 U17877 ( .B(n25487), .A(n25494), .S(n27711), .Y(n27409) );
  MUX2X1 U17878 ( .B(n27408), .A(n27405), .S(n27702), .Y(n27419) );
  MUX2X1 U17879 ( .B(grid[229]), .A(grid[235]), .S(n27711), .Y(n27413) );
  MUX2X1 U17880 ( .B(grid[217]), .A(n20831), .S(n27711), .Y(n27412) );
  MUX2X1 U17881 ( .B(n25600), .A(n25481), .S(n27711), .Y(n27416) );
  MUX2X1 U17882 ( .B(grid[193]), .A(grid[199]), .S(n27711), .Y(n27415) );
  MUX2X1 U17883 ( .B(n27414), .A(n27411), .S(n27702), .Y(n27418) );
  MUX2X1 U17884 ( .B(n27417), .A(n27402), .S(n20812), .Y(n27451) );
  MUX2X1 U17885 ( .B(grid[181]), .A(n25496), .S(n27710), .Y(n27422) );
  MUX2X1 U17886 ( .B(grid[169]), .A(grid[175]), .S(n27710), .Y(n27421) );
  MUX2X1 U17887 ( .B(grid[157]), .A(grid[163]), .S(n27710), .Y(n27425) );
  MUX2X1 U17888 ( .B(grid[145]), .A(grid[151]), .S(n27710), .Y(n27424) );
  MUX2X1 U17889 ( .B(n27423), .A(n27420), .S(n27702), .Y(n27434) );
  MUX2X1 U17890 ( .B(grid[133]), .A(grid[139]), .S(n27710), .Y(n27428) );
  MUX2X1 U17891 ( .B(grid[121]), .A(grid[127]), .S(n27710), .Y(n27427) );
  MUX2X1 U17892 ( .B(grid[109]), .A(grid[115]), .S(n27710), .Y(n27431) );
  MUX2X1 U17893 ( .B(grid[97]), .A(n25516), .S(n27710), .Y(n27430) );
  MUX2X1 U17894 ( .B(n27429), .A(n27426), .S(n27702), .Y(n27433) );
  MUX2X1 U17895 ( .B(grid[85]), .A(n25501), .S(n27710), .Y(n27437) );
  MUX2X1 U17896 ( .B(n25578), .A(grid[79]), .S(n27710), .Y(n27436) );
  MUX2X1 U17897 ( .B(n25622), .A(grid[67]), .S(n27710), .Y(n27440) );
  MUX2X1 U17898 ( .B(n25607), .A(n25512), .S(n27710), .Y(n27439) );
  MUX2X1 U17899 ( .B(n27438), .A(n27435), .S(n27702), .Y(n27449) );
  MUX2X1 U17900 ( .B(n25608), .A(n25577), .S(n27709), .Y(n27443) );
  MUX2X1 U17901 ( .B(grid[25]), .A(n25603), .S(n27709), .Y(n27442) );
  MUX2X1 U17902 ( .B(grid[13]), .A(grid[19]), .S(n27709), .Y(n27446) );
  MUX2X1 U17903 ( .B(grid[1]), .A(grid[7]), .S(n27709), .Y(n27445) );
  MUX2X1 U17904 ( .B(n27444), .A(n27441), .S(n27702), .Y(n27448) );
  MUX2X1 U17905 ( .B(n27447), .A(n27432), .S(n20812), .Y(n27450) );
  MUX2X1 U17906 ( .B(grid[374]), .A(grid[380]), .S(n27709), .Y(n27454) );
  MUX2X1 U17907 ( .B(grid[362]), .A(grid[368]), .S(n27709), .Y(n27453) );
  MUX2X1 U17908 ( .B(grid[350]), .A(grid[356]), .S(n27709), .Y(n27457) );
  MUX2X1 U17909 ( .B(n25500), .A(grid[344]), .S(n27709), .Y(n27456) );
  MUX2X1 U17910 ( .B(n27455), .A(n27452), .S(n27702), .Y(n27466) );
  MUX2X1 U17911 ( .B(n25502), .A(grid[332]), .S(n27709), .Y(n27460) );
  MUX2X1 U17912 ( .B(grid[314]), .A(grid[320]), .S(n27709), .Y(n27459) );
  MUX2X1 U17913 ( .B(n25605), .A(grid[308]), .S(n27709), .Y(n27463) );
  MUX2X1 U17914 ( .B(n25610), .A(grid[296]), .S(n27709), .Y(n27462) );
  MUX2X1 U17915 ( .B(n27461), .A(n27458), .S(n27702), .Y(n27465) );
  MUX2X1 U17916 ( .B(n25465), .A(grid[284]), .S(n27708), .Y(n27469) );
  MUX2X1 U17917 ( .B(n25598), .A(grid[272]), .S(n27708), .Y(n27468) );
  MUX2X1 U17918 ( .B(grid[254]), .A(n25602), .S(n27708), .Y(n27472) );
  MUX2X1 U17919 ( .B(n25660), .A(grid[248]), .S(n27708), .Y(n27471) );
  MUX2X1 U17920 ( .B(n27470), .A(n27467), .S(n27702), .Y(n27481) );
  MUX2X1 U17921 ( .B(n25509), .A(grid[236]), .S(n27708), .Y(n27475) );
  MUX2X1 U17922 ( .B(grid[218]), .A(grid[224]), .S(n27708), .Y(n27474) );
  MUX2X1 U17923 ( .B(n25654), .A(grid[212]), .S(n27708), .Y(n27478) );
  MUX2X1 U17924 ( .B(n25599), .A(n25514), .S(n27708), .Y(n27477) );
  MUX2X1 U17925 ( .B(n27476), .A(n27473), .S(n27702), .Y(n27480) );
  MUX2X1 U17926 ( .B(n27479), .A(n27464), .S(n20812), .Y(n27513) );
  MUX2X1 U17927 ( .B(grid[182]), .A(grid[188]), .S(n27708), .Y(n27484) );
  MUX2X1 U17928 ( .B(grid[170]), .A(grid[176]), .S(n27708), .Y(n27483) );
  MUX2X1 U17929 ( .B(n25595), .A(grid[164]), .S(n27708), .Y(n27487) );
  MUX2X1 U17930 ( .B(n25574), .A(grid[152]), .S(n27708), .Y(n27486) );
  MUX2X1 U17931 ( .B(n27485), .A(n27482), .S(n27702), .Y(n27496) );
  MUX2X1 U17932 ( .B(grid[134]), .A(grid[140]), .S(n27707), .Y(n27490) );
  MUX2X1 U17933 ( .B(grid[122]), .A(grid[128]), .S(n27707), .Y(n27489) );
  MUX2X1 U17934 ( .B(n25601), .A(grid[116]), .S(n27707), .Y(n27493) );
  MUX2X1 U17935 ( .B(n25495), .A(grid[104]), .S(n27707), .Y(n27492) );
  MUX2X1 U17936 ( .B(n27491), .A(n27488), .S(n27702), .Y(n27495) );
  MUX2X1 U17937 ( .B(grid[86]), .A(grid[92]), .S(n27707), .Y(n27499) );
  MUX2X1 U17938 ( .B(n25503), .A(grid[80]), .S(n27707), .Y(n27498) );
  MUX2X1 U17939 ( .B(n25659), .A(grid[68]), .S(n27707), .Y(n27502) );
  MUX2X1 U17940 ( .B(n25655), .A(n25581), .S(n27707), .Y(n27501) );
  MUX2X1 U17941 ( .B(n27500), .A(n27497), .S(n27702), .Y(n27511) );
  MUX2X1 U17942 ( .B(n25508), .A(grid[44]), .S(n27707), .Y(n27505) );
  MUX2X1 U17943 ( .B(n25484), .A(grid[32]), .S(n27707), .Y(n27504) );
  MUX2X1 U17944 ( .B(n25656), .A(n25582), .S(n27707), .Y(n27508) );
  MUX2X1 U17945 ( .B(n25576), .A(grid[8]), .S(n27707), .Y(n27507) );
  MUX2X1 U17946 ( .B(n27506), .A(n27503), .S(n27702), .Y(n27510) );
  MUX2X1 U17947 ( .B(n27509), .A(n27494), .S(n20812), .Y(n27512) );
  MUX2X1 U17948 ( .B(grid[375]), .A(grid[381]), .S(n27706), .Y(n27516) );
  MUX2X1 U17949 ( .B(grid[363]), .A(grid[369]), .S(n27706), .Y(n27515) );
  MUX2X1 U17950 ( .B(grid[351]), .A(grid[357]), .S(n27706), .Y(n27519) );
  MUX2X1 U17951 ( .B(grid[339]), .A(grid[345]), .S(n27706), .Y(n27518) );
  MUX2X1 U17952 ( .B(n27517), .A(n27514), .S(n27702), .Y(n27528) );
  MUX2X1 U17953 ( .B(grid[327]), .A(grid[333]), .S(n27706), .Y(n27522) );
  MUX2X1 U17954 ( .B(grid[315]), .A(grid[321]), .S(n27706), .Y(n27521) );
  MUX2X1 U17955 ( .B(grid[303]), .A(grid[309]), .S(n27706), .Y(n27525) );
  MUX2X1 U17956 ( .B(grid[291]), .A(grid[297]), .S(n27706), .Y(n27524) );
  MUX2X1 U17957 ( .B(n27523), .A(n27520), .S(n27702), .Y(n27527) );
  MUX2X1 U17958 ( .B(grid[279]), .A(grid[285]), .S(n27706), .Y(n27531) );
  MUX2X1 U17959 ( .B(grid[267]), .A(grid[273]), .S(n27706), .Y(n27530) );
  MUX2X1 U17960 ( .B(grid[255]), .A(grid[261]), .S(n27706), .Y(n27534) );
  MUX2X1 U17961 ( .B(grid[243]), .A(grid[249]), .S(n27706), .Y(n27533) );
  MUX2X1 U17962 ( .B(n27532), .A(n27529), .S(n27702), .Y(n27543) );
  MUX2X1 U17963 ( .B(grid[231]), .A(grid[237]), .S(n27705), .Y(n27537) );
  MUX2X1 U17964 ( .B(grid[219]), .A(grid[225]), .S(n27705), .Y(n27536) );
  MUX2X1 U17965 ( .B(grid[207]), .A(grid[213]), .S(n27705), .Y(n27540) );
  MUX2X1 U17966 ( .B(grid[195]), .A(grid[201]), .S(n27705), .Y(n27539) );
  MUX2X1 U17967 ( .B(n27538), .A(n27535), .S(n27702), .Y(n27542) );
  MUX2X1 U17968 ( .B(n27541), .A(n27526), .S(n20812), .Y(n27575) );
  MUX2X1 U17969 ( .B(grid[183]), .A(grid[189]), .S(n27705), .Y(n27546) );
  MUX2X1 U17970 ( .B(grid[171]), .A(grid[177]), .S(n27705), .Y(n27545) );
  MUX2X1 U17971 ( .B(grid[159]), .A(grid[165]), .S(n27705), .Y(n27549) );
  MUX2X1 U17972 ( .B(grid[147]), .A(grid[153]), .S(n27705), .Y(n27548) );
  MUX2X1 U17973 ( .B(n27547), .A(n27544), .S(n27702), .Y(n27558) );
  MUX2X1 U17974 ( .B(grid[135]), .A(grid[141]), .S(n27705), .Y(n27552) );
  MUX2X1 U17975 ( .B(grid[123]), .A(grid[129]), .S(n27705), .Y(n27551) );
  MUX2X1 U17976 ( .B(grid[111]), .A(grid[117]), .S(n27705), .Y(n27555) );
  MUX2X1 U17977 ( .B(grid[99]), .A(grid[105]), .S(n27705), .Y(n27554) );
  MUX2X1 U17978 ( .B(n27553), .A(n27550), .S(n27702), .Y(n27557) );
  MUX2X1 U17979 ( .B(grid[87]), .A(grid[93]), .S(n27711), .Y(n27561) );
  MUX2X1 U17980 ( .B(grid[75]), .A(grid[81]), .S(n27707), .Y(n27560) );
  MUX2X1 U17981 ( .B(grid[63]), .A(grid[69]), .S(n27713), .Y(n27564) );
  MUX2X1 U17982 ( .B(grid[51]), .A(grid[57]), .S(n27705), .Y(n27563) );
  MUX2X1 U17983 ( .B(n27562), .A(n27559), .S(n27702), .Y(n27573) );
  MUX2X1 U17984 ( .B(grid[39]), .A(grid[45]), .S(n27708), .Y(n27567) );
  MUX2X1 U17985 ( .B(grid[27]), .A(grid[33]), .S(n27712), .Y(n27566) );
  MUX2X1 U17986 ( .B(grid[15]), .A(grid[21]), .S(n27714), .Y(n27570) );
  MUX2X1 U17987 ( .B(grid[3]), .A(grid[9]), .S(n27706), .Y(n27569) );
  MUX2X1 U17988 ( .B(n27568), .A(n27565), .S(n27702), .Y(n27572) );
  MUX2X1 U17989 ( .B(n27571), .A(n27556), .S(n20812), .Y(n27574) );
  MUX2X1 U17990 ( .B(grid[376]), .A(grid[382]), .S(n20978), .Y(n27578) );
  MUX2X1 U17991 ( .B(grid[364]), .A(grid[370]), .S(n27709), .Y(n27577) );
  MUX2X1 U17992 ( .B(grid[352]), .A(grid[358]), .S(n27710), .Y(n27581) );
  MUX2X1 U17993 ( .B(grid[340]), .A(grid[346]), .S(n27711), .Y(n27580) );
  MUX2X1 U17994 ( .B(n27579), .A(n27576), .S(n27702), .Y(n27590) );
  MUX2X1 U17995 ( .B(grid[328]), .A(grid[334]), .S(n27712), .Y(n27584) );
  MUX2X1 U17996 ( .B(grid[316]), .A(grid[322]), .S(n27714), .Y(n27583) );
  MUX2X1 U17997 ( .B(grid[304]), .A(grid[310]), .S(n27706), .Y(n27587) );
  MUX2X1 U17998 ( .B(grid[292]), .A(grid[298]), .S(n20978), .Y(n27586) );
  MUX2X1 U17999 ( .B(n27585), .A(n27582), .S(n27702), .Y(n27589) );
  MUX2X1 U18000 ( .B(grid[280]), .A(grid[286]), .S(n27709), .Y(n27593) );
  MUX2X1 U18001 ( .B(grid[268]), .A(grid[274]), .S(n27710), .Y(n27592) );
  MUX2X1 U18002 ( .B(grid[256]), .A(grid[262]), .S(n27711), .Y(n27596) );
  MUX2X1 U18003 ( .B(grid[244]), .A(grid[250]), .S(n27707), .Y(n27595) );
  MUX2X1 U18004 ( .B(n27594), .A(n27591), .S(n27702), .Y(n27605) );
  MUX2X1 U18005 ( .B(grid[232]), .A(grid[238]), .S(n27708), .Y(n27599) );
  MUX2X1 U18006 ( .B(grid[220]), .A(grid[226]), .S(n27713), .Y(n27598) );
  MUX2X1 U18007 ( .B(grid[208]), .A(grid[214]), .S(n27705), .Y(n27602) );
  MUX2X1 U18008 ( .B(grid[196]), .A(grid[202]), .S(n27708), .Y(n27601) );
  MUX2X1 U18009 ( .B(n27600), .A(n27597), .S(n27702), .Y(n27604) );
  MUX2X1 U18010 ( .B(n27603), .A(n27588), .S(n20812), .Y(n27637) );
  MUX2X1 U18011 ( .B(grid[184]), .A(grid[190]), .S(n20978), .Y(n27608) );
  MUX2X1 U18012 ( .B(grid[172]), .A(grid[178]), .S(n27709), .Y(n27607) );
  MUX2X1 U18013 ( .B(grid[160]), .A(grid[166]), .S(n27710), .Y(n27611) );
  MUX2X1 U18014 ( .B(grid[148]), .A(grid[154]), .S(n27711), .Y(n27610) );
  MUX2X1 U18015 ( .B(n27609), .A(n27606), .S(n27702), .Y(n27620) );
  MUX2X1 U18016 ( .B(grid[136]), .A(grid[142]), .S(n27707), .Y(n27614) );
  MUX2X1 U18017 ( .B(grid[124]), .A(grid[130]), .S(n27705), .Y(n27613) );
  MUX2X1 U18018 ( .B(grid[112]), .A(grid[118]), .S(n27713), .Y(n27617) );
  MUX2X1 U18019 ( .B(grid[100]), .A(grid[106]), .S(n27705), .Y(n27616) );
  MUX2X1 U18020 ( .B(n27615), .A(n27612), .S(n27702), .Y(n27619) );
  MUX2X1 U18021 ( .B(grid[88]), .A(grid[94]), .S(n27706), .Y(n27623) );
  MUX2X1 U18022 ( .B(grid[76]), .A(grid[82]), .S(n27708), .Y(n27622) );
  MUX2X1 U18023 ( .B(grid[64]), .A(grid[70]), .S(n27712), .Y(n27626) );
  MUX2X1 U18024 ( .B(grid[52]), .A(grid[58]), .S(n27714), .Y(n27625) );
  MUX2X1 U18025 ( .B(n27624), .A(n27621), .S(n27702), .Y(n27635) );
  MUX2X1 U18026 ( .B(grid[40]), .A(grid[46]), .S(n27709), .Y(n27629) );
  MUX2X1 U18027 ( .B(grid[28]), .A(grid[34]), .S(n27710), .Y(n27628) );
  MUX2X1 U18028 ( .B(grid[16]), .A(grid[22]), .S(n27711), .Y(n27632) );
  MUX2X1 U18029 ( .B(grid[4]), .A(grid[10]), .S(n27707), .Y(n27631) );
  MUX2X1 U18030 ( .B(n27630), .A(n27627), .S(n27702), .Y(n27634) );
  MUX2X1 U18031 ( .B(n27633), .A(n27618), .S(n20812), .Y(n27636) );
  MUX2X1 U18032 ( .B(grid[377]), .A(grid[383]), .S(n27713), .Y(n27640) );
  MUX2X1 U18033 ( .B(grid[365]), .A(grid[371]), .S(n27713), .Y(n27639) );
  MUX2X1 U18034 ( .B(grid[353]), .A(grid[359]), .S(n27705), .Y(n27643) );
  MUX2X1 U18035 ( .B(grid[341]), .A(grid[347]), .S(n20978), .Y(n27642) );
  MUX2X1 U18036 ( .B(n27641), .A(n27638), .S(n27702), .Y(n27652) );
  MUX2X1 U18037 ( .B(grid[329]), .A(grid[335]), .S(n27714), .Y(n27646) );
  MUX2X1 U18038 ( .B(grid[317]), .A(grid[323]), .S(n27708), .Y(n27645) );
  MUX2X1 U18039 ( .B(grid[305]), .A(grid[311]), .S(n27712), .Y(n27649) );
  MUX2X1 U18040 ( .B(grid[293]), .A(grid[299]), .S(n27714), .Y(n27648) );
  MUX2X1 U18041 ( .B(n27647), .A(n27644), .S(n27702), .Y(n27651) );
  MUX2X1 U18042 ( .B(grid[281]), .A(grid[287]), .S(n20978), .Y(n27655) );
  MUX2X1 U18043 ( .B(grid[269]), .A(grid[275]), .S(n27709), .Y(n27654) );
  MUX2X1 U18044 ( .B(grid[257]), .A(grid[263]), .S(n27710), .Y(n27658) );
  MUX2X1 U18045 ( .B(grid[245]), .A(grid[251]), .S(n27711), .Y(n27657) );
  MUX2X1 U18046 ( .B(n27656), .A(n27653), .S(n27702), .Y(n27667) );
  MUX2X1 U18047 ( .B(grid[233]), .A(grid[239]), .S(n27707), .Y(n27661) );
  MUX2X1 U18048 ( .B(grid[221]), .A(grid[227]), .S(n27707), .Y(n27660) );
  MUX2X1 U18049 ( .B(grid[209]), .A(grid[215]), .S(n27713), .Y(n27664) );
  MUX2X1 U18050 ( .B(grid[197]), .A(grid[203]), .S(n27705), .Y(n27663) );
  MUX2X1 U18051 ( .B(n27662), .A(n27659), .S(n27702), .Y(n27666) );
  MUX2X1 U18052 ( .B(n27665), .A(n27650), .S(n20812), .Y(n27699) );
  MUX2X1 U18053 ( .B(grid[185]), .A(grid[191]), .S(n27706), .Y(n27670) );
  MUX2X1 U18054 ( .B(grid[173]), .A(grid[179]), .S(n27706), .Y(n27669) );
  MUX2X1 U18055 ( .B(grid[161]), .A(grid[167]), .S(n27712), .Y(n27673) );
  MUX2X1 U18056 ( .B(grid[149]), .A(grid[155]), .S(n27708), .Y(n27672) );
  MUX2X1 U18057 ( .B(n27671), .A(n27668), .S(n27702), .Y(n27682) );
  MUX2X1 U18058 ( .B(grid[137]), .A(grid[143]), .S(n27712), .Y(n27676) );
  MUX2X1 U18059 ( .B(grid[125]), .A(grid[131]), .S(n27714), .Y(n27675) );
  MUX2X1 U18060 ( .B(grid[113]), .A(grid[119]), .S(n27706), .Y(n27679) );
  MUX2X1 U18061 ( .B(grid[101]), .A(grid[107]), .S(n20978), .Y(n27678) );
  MUX2X1 U18062 ( .B(n27677), .A(n27674), .S(n27702), .Y(n27681) );
  MUX2X1 U18063 ( .B(grid[89]), .A(grid[95]), .S(n20978), .Y(n27685) );
  MUX2X1 U18064 ( .B(grid[77]), .A(grid[83]), .S(n20978), .Y(n27684) );
  MUX2X1 U18065 ( .B(grid[65]), .A(grid[71]), .S(n20978), .Y(n27688) );
  MUX2X1 U18066 ( .B(grid[53]), .A(grid[59]), .S(n20978), .Y(n27687) );
  MUX2X1 U18067 ( .B(n27686), .A(n27683), .S(n27702), .Y(n27697) );
  MUX2X1 U18068 ( .B(grid[41]), .A(grid[47]), .S(n20978), .Y(n27691) );
  MUX2X1 U18069 ( .B(grid[29]), .A(grid[35]), .S(n20978), .Y(n27690) );
  MUX2X1 U18070 ( .B(grid[17]), .A(grid[23]), .S(n20978), .Y(n27694) );
  MUX2X1 U18071 ( .B(grid[5]), .A(grid[11]), .S(n20978), .Y(n27693) );
  MUX2X1 U18072 ( .B(n27692), .A(n27689), .S(n27702), .Y(n27696) );
  MUX2X1 U18073 ( .B(n27695), .A(n27680), .S(n20812), .Y(n27698) );
  MUX2X1 U18074 ( .B(n27717), .A(n27718), .S(n27911), .Y(n27716) );
  MUX2X1 U18075 ( .B(n27720), .A(n27721), .S(n27911), .Y(n27719) );
  MUX2X1 U18076 ( .B(n27723), .A(n27724), .S(n27912), .Y(n27722) );
  MUX2X1 U18077 ( .B(n27726), .A(n27727), .S(n27911), .Y(n27725) );
  MUX2X1 U18078 ( .B(n27729), .A(n27730), .S(n25620), .Y(n27728) );
  MUX2X1 U18079 ( .B(n27732), .A(n27733), .S(n27911), .Y(n27731) );
  MUX2X1 U18080 ( .B(n27735), .A(n27736), .S(n27911), .Y(n27734) );
  MUX2X1 U18081 ( .B(n27738), .A(n27739), .S(n27912), .Y(n27737) );
  MUX2X1 U18082 ( .B(n27741), .A(n27742), .S(n27911), .Y(n27740) );
  MUX2X1 U18083 ( .B(n27744), .A(n27745), .S(n27917), .Y(n27743) );
  MUX2X1 U18084 ( .B(n27747), .A(n27748), .S(n27911), .Y(n27746) );
  MUX2X1 U18085 ( .B(n27750), .A(n27751), .S(n27911), .Y(n27749) );
  MUX2X1 U18086 ( .B(n27753), .A(n27754), .S(n27911), .Y(n27752) );
  MUX2X1 U18087 ( .B(n27756), .A(n27757), .S(n27912), .Y(n27755) );
  MUX2X1 U18088 ( .B(n27759), .A(n27760), .S(n27916), .Y(n27758) );
  MUX2X1 U18089 ( .B(n27762), .A(n27763), .S(n27911), .Y(n27761) );
  MUX2X1 U18090 ( .B(n27765), .A(n27766), .S(n27911), .Y(n27764) );
  MUX2X1 U18091 ( .B(n27768), .A(n27769), .S(n27911), .Y(n27767) );
  MUX2X1 U18092 ( .B(n27771), .A(n27772), .S(n27911), .Y(n27770) );
  MUX2X1 U18093 ( .B(n27774), .A(n27775), .S(n25649), .Y(n27773) );
  MUX2X1 U18094 ( .B(n27776), .A(n27777), .S(n20969), .Y(n3774) );
  MUX2X1 U18095 ( .B(n27779), .A(n27780), .S(n27911), .Y(n27778) );
  MUX2X1 U18096 ( .B(n27782), .A(n27783), .S(n27911), .Y(n27781) );
  MUX2X1 U18097 ( .B(n27785), .A(n27786), .S(n27911), .Y(n27784) );
  MUX2X1 U18098 ( .B(n27788), .A(n27789), .S(n27911), .Y(n27787) );
  MUX2X1 U18099 ( .B(n27794), .A(n27795), .S(n27911), .Y(n27793) );
  MUX2X1 U18100 ( .B(n27797), .A(n27798), .S(n27911), .Y(n27796) );
  MUX2X1 U18101 ( .B(n27800), .A(n27801), .S(n27911), .Y(n27799) );
  MUX2X1 U18102 ( .B(n27803), .A(n27804), .S(n27911), .Y(n27802) );
  MUX2X1 U18103 ( .B(n27806), .A(n27807), .S(n25621), .Y(n27805) );
  MUX2X1 U18104 ( .B(n27809), .A(n27810), .S(n27911), .Y(n27808) );
  MUX2X1 U18105 ( .B(n27812), .A(n27813), .S(n27911), .Y(n27811) );
  MUX2X1 U18106 ( .B(n27815), .A(n27816), .S(n27912), .Y(n27814) );
  MUX2X1 U18107 ( .B(n27818), .A(n27819), .S(n27911), .Y(n27817) );
  MUX2X1 U18108 ( .B(n27821), .A(n27822), .S(n25620), .Y(n27820) );
  MUX2X1 U18109 ( .B(n27824), .A(n27825), .S(n27911), .Y(n27823) );
  MUX2X1 U18110 ( .B(n27827), .A(n27828), .S(n27911), .Y(n27826) );
  MUX2X1 U18111 ( .B(n27830), .A(n27831), .S(n27911), .Y(n27829) );
  MUX2X1 U18112 ( .B(n27833), .A(n27834), .S(n27912), .Y(n27832) );
  MUX2X1 U18113 ( .B(n27836), .A(n27837), .S(n25621), .Y(n27835) );
  MUX2X1 U18114 ( .B(n27838), .A(n27839), .S(n20969), .Y(n3773) );
  MUX2X1 U18115 ( .B(n27841), .A(n27842), .S(n27911), .Y(n27840) );
  MUX2X1 U18116 ( .B(n27844), .A(n27845), .S(n27911), .Y(n27843) );
  MUX2X1 U18117 ( .B(n27847), .A(n27848), .S(n27911), .Y(n27846) );
  MUX2X1 U18118 ( .B(n27850), .A(n27851), .S(n27911), .Y(n27849) );
  MUX2X1 U18119 ( .B(n27853), .A(n27854), .S(n25649), .Y(n27852) );
  MUX2X1 U18120 ( .B(n27856), .A(n27857), .S(n27911), .Y(n27855) );
  MUX2X1 U18121 ( .B(n27859), .A(n27860), .S(n27911), .Y(n27858) );
  MUX2X1 U18122 ( .B(n27862), .A(n27863), .S(n27911), .Y(n27861) );
  MUX2X1 U18123 ( .B(n27865), .A(n27866), .S(n27911), .Y(n27864) );
  MUX2X1 U18124 ( .B(n27868), .A(n27869), .S(n25649), .Y(n27867) );
  MUX2X1 U18125 ( .B(n27871), .A(n27872), .S(n27911), .Y(n27870) );
  MUX2X1 U18126 ( .B(n27874), .A(n27875), .S(n27911), .Y(n27873) );
  MUX2X1 U18127 ( .B(n27877), .A(n27878), .S(n27911), .Y(n27876) );
  MUX2X1 U18128 ( .B(n27880), .A(n27881), .S(n27911), .Y(n27879) );
  MUX2X1 U18129 ( .B(n27883), .A(n27884), .S(n25621), .Y(n27882) );
  MUX2X1 U18130 ( .B(n27886), .A(n27887), .S(n27912), .Y(n27885) );
  MUX2X1 U18131 ( .B(n27889), .A(n27890), .S(n27911), .Y(n27888) );
  MUX2X1 U18132 ( .B(n27892), .A(n27893), .S(n27911), .Y(n27891) );
  MUX2X1 U18133 ( .B(n27895), .A(n27896), .S(n27911), .Y(n27894) );
  MUX2X1 U18134 ( .B(n27898), .A(n27899), .S(n25620), .Y(n27897) );
  MUX2X1 U18135 ( .B(n27900), .A(n27901), .S(n20969), .Y(n3772) );
  MUX2X1 U18136 ( .B(grid[372]), .A(grid[378]), .S(n27910), .Y(n27718) );
  MUX2X1 U18137 ( .B(n21081), .A(grid[366]), .S(n27910), .Y(n27717) );
  MUX2X1 U18138 ( .B(n25626), .A(grid[354]), .S(n27910), .Y(n27721) );
  MUX2X1 U18139 ( .B(grid[336]), .A(grid[342]), .S(n27910), .Y(n27720) );
  MUX2X1 U18140 ( .B(n27719), .A(n27716), .S(n27914), .Y(n27730) );
  MUX2X1 U18141 ( .B(grid[324]), .A(grid[330]), .S(n27910), .Y(n27724) );
  MUX2X1 U18142 ( .B(grid[312]), .A(grid[318]), .S(n27910), .Y(n27723) );
  MUX2X1 U18143 ( .B(n25618), .A(grid[306]), .S(n27910), .Y(n27727) );
  MUX2X1 U18144 ( .B(grid[288]), .A(grid[294]), .S(n27910), .Y(n27726) );
  MUX2X1 U18145 ( .B(n27725), .A(n27722), .S(n27914), .Y(n27729) );
  MUX2X1 U18146 ( .B(n25627), .A(grid[282]), .S(n27910), .Y(n27733) );
  MUX2X1 U18147 ( .B(grid[264]), .A(grid[270]), .S(n27910), .Y(n27732) );
  MUX2X1 U18148 ( .B(n25643), .A(grid[258]), .S(n27910), .Y(n27736) );
  MUX2X1 U18149 ( .B(n25637), .A(grid[246]), .S(n27910), .Y(n27735) );
  MUX2X1 U18150 ( .B(n27734), .A(n27731), .S(n27914), .Y(n27745) );
  MUX2X1 U18151 ( .B(n21088), .A(grid[234]), .S(n27909), .Y(n27739) );
  MUX2X1 U18152 ( .B(grid[216]), .A(grid[222]), .S(n27909), .Y(n27738) );
  MUX2X1 U18153 ( .B(n25635), .A(grid[210]), .S(n27909), .Y(n27742) );
  MUX2X1 U18154 ( .B(n25631), .A(grid[198]), .S(n27909), .Y(n27741) );
  MUX2X1 U18155 ( .B(n27740), .A(n27737), .S(n27914), .Y(n27744) );
  MUX2X1 U18156 ( .B(n27743), .A(n27728), .S(n25619), .Y(n27777) );
  MUX2X1 U18157 ( .B(grid[180]), .A(grid[186]), .S(n20850), .Y(n27748) );
  MUX2X1 U18158 ( .B(grid[168]), .A(grid[174]), .S(n20850), .Y(n27747) );
  MUX2X1 U18159 ( .B(grid[156]), .A(n25625), .S(n27909), .Y(n27751) );
  MUX2X1 U18160 ( .B(n21084), .A(grid[150]), .S(n27909), .Y(n27750) );
  MUX2X1 U18161 ( .B(n27749), .A(n27746), .S(n27914), .Y(n27760) );
  MUX2X1 U18162 ( .B(grid[132]), .A(grid[138]), .S(n20850), .Y(n27754) );
  MUX2X1 U18163 ( .B(grid[120]), .A(grid[126]), .S(n20850), .Y(n27753) );
  MUX2X1 U18164 ( .B(grid[108]), .A(grid[114]), .S(n27909), .Y(n27757) );
  MUX2X1 U18165 ( .B(grid[96]), .A(grid[102]), .S(n20850), .Y(n27756) );
  MUX2X1 U18166 ( .B(n27755), .A(n27752), .S(n27914), .Y(n27759) );
  MUX2X1 U18167 ( .B(grid[84]), .A(n21082), .S(n25685), .Y(n27763) );
  MUX2X1 U18168 ( .B(grid[72]), .A(grid[78]), .S(n27909), .Y(n27762) );
  MUX2X1 U18169 ( .B(n25639), .A(grid[66]), .S(n27907), .Y(n27766) );
  MUX2X1 U18170 ( .B(n25632), .A(grid[54]), .S(n25685), .Y(n27765) );
  MUX2X1 U18171 ( .B(n27764), .A(n27761), .S(n27914), .Y(n27775) );
  MUX2X1 U18172 ( .B(n21087), .A(grid[42]), .S(n27909), .Y(n27769) );
  MUX2X1 U18173 ( .B(grid[24]), .A(grid[30]), .S(n20850), .Y(n27768) );
  MUX2X1 U18174 ( .B(n25633), .A(grid[18]), .S(n25685), .Y(n27772) );
  MUX2X1 U18175 ( .B(grid[0]), .A(n21086), .S(n27909), .Y(n27771) );
  MUX2X1 U18176 ( .B(n27770), .A(n27767), .S(n27914), .Y(n27774) );
  MUX2X1 U18177 ( .B(n27773), .A(n27758), .S(n25688), .Y(n27776) );
  MUX2X1 U18178 ( .B(grid[373]), .A(grid[379]), .S(n27909), .Y(n27780) );
  MUX2X1 U18179 ( .B(grid[349]), .A(n25486), .S(n27909), .Y(n27783) );
  MUX2X1 U18180 ( .B(grid[337]), .A(n25492), .S(n27909), .Y(n27782) );
  MUX2X1 U18181 ( .B(n27781), .A(n27778), .S(n27914), .Y(n27792) );
  MUX2X1 U18182 ( .B(grid[325]), .A(n23205), .S(n27907), .Y(n27786) );
  MUX2X1 U18183 ( .B(grid[313]), .A(grid[319]), .S(n27910), .Y(n27785) );
  MUX2X1 U18184 ( .B(n20845), .A(n25493), .S(n27907), .Y(n27789) );
  MUX2X1 U18185 ( .B(grid[289]), .A(grid[295]), .S(n25711), .Y(n27788) );
  MUX2X1 U18186 ( .B(n27787), .A(n27784), .S(n27914), .Y(n27791) );
  MUX2X1 U18187 ( .B(n25513), .A(grid[283]), .S(n27907), .Y(n27795) );
  MUX2X1 U18188 ( .B(n25506), .A(grid[271]), .S(n27907), .Y(n27794) );
  MUX2X1 U18189 ( .B(n25490), .A(grid[259]), .S(n25685), .Y(n27798) );
  MUX2X1 U18190 ( .B(n25487), .A(n25494), .S(n25711), .Y(n27797) );
  MUX2X1 U18191 ( .B(n27796), .A(n27793), .S(n27914), .Y(n27807) );
  MUX2X1 U18192 ( .B(grid[229]), .A(grid[235]), .S(n25685), .Y(n27801) );
  MUX2X1 U18193 ( .B(grid[217]), .A(n20831), .S(n25685), .Y(n27800) );
  MUX2X1 U18194 ( .B(n25600), .A(grid[211]), .S(n25685), .Y(n27804) );
  MUX2X1 U18195 ( .B(grid[193]), .A(grid[199]), .S(n25685), .Y(n27803) );
  MUX2X1 U18196 ( .B(n27802), .A(n27799), .S(n27914), .Y(n27806) );
  MUX2X1 U18197 ( .B(n27805), .A(n27790), .S(n25619), .Y(n27839) );
  MUX2X1 U18198 ( .B(grid[181]), .A(n25496), .S(n27908), .Y(n27810) );
  MUX2X1 U18199 ( .B(grid[169]), .A(grid[175]), .S(n27908), .Y(n27809) );
  MUX2X1 U18200 ( .B(grid[157]), .A(grid[163]), .S(n27908), .Y(n27813) );
  MUX2X1 U18201 ( .B(grid[145]), .A(grid[151]), .S(n27908), .Y(n27812) );
  MUX2X1 U18202 ( .B(n27811), .A(n27808), .S(n27914), .Y(n27822) );
  MUX2X1 U18203 ( .B(grid[133]), .A(grid[139]), .S(n27908), .Y(n27816) );
  MUX2X1 U18204 ( .B(grid[121]), .A(grid[127]), .S(n27908), .Y(n27815) );
  MUX2X1 U18205 ( .B(grid[109]), .A(grid[115]), .S(n27908), .Y(n27819) );
  MUX2X1 U18206 ( .B(grid[97]), .A(n25516), .S(n27908), .Y(n27818) );
  MUX2X1 U18207 ( .B(n27817), .A(n27814), .S(n27914), .Y(n27821) );
  MUX2X1 U18208 ( .B(grid[85]), .A(n25501), .S(n27908), .Y(n27825) );
  MUX2X1 U18209 ( .B(n25578), .A(grid[79]), .S(n27908), .Y(n27824) );
  MUX2X1 U18210 ( .B(n25622), .A(grid[67]), .S(n27908), .Y(n27828) );
  MUX2X1 U18211 ( .B(n25607), .A(n25497), .S(n27908), .Y(n27827) );
  MUX2X1 U18212 ( .B(n27826), .A(n27823), .S(n27914), .Y(n27837) );
  MUX2X1 U18213 ( .B(n25608), .A(n25507), .S(n25685), .Y(n27831) );
  MUX2X1 U18214 ( .B(grid[25]), .A(grid[31]), .S(n27907), .Y(n27830) );
  MUX2X1 U18215 ( .B(grid[13]), .A(grid[19]), .S(n25711), .Y(n27834) );
  MUX2X1 U18216 ( .B(grid[1]), .A(grid[7]), .S(n25711), .Y(n27833) );
  MUX2X1 U18217 ( .B(n27832), .A(n27829), .S(n27914), .Y(n27836) );
  MUX2X1 U18218 ( .B(n27835), .A(n27820), .S(n25688), .Y(n27838) );
  MUX2X1 U18219 ( .B(grid[374]), .A(grid[380]), .S(n27907), .Y(n27842) );
  MUX2X1 U18220 ( .B(grid[362]), .A(grid[368]), .S(n25711), .Y(n27841) );
  MUX2X1 U18221 ( .B(grid[350]), .A(grid[356]), .S(n25711), .Y(n27845) );
  MUX2X1 U18222 ( .B(n25500), .A(grid[344]), .S(n27907), .Y(n27844) );
  MUX2X1 U18223 ( .B(n27843), .A(n27840), .S(n27914), .Y(n27854) );
  MUX2X1 U18224 ( .B(n25502), .A(grid[332]), .S(n25711), .Y(n27848) );
  MUX2X1 U18225 ( .B(grid[314]), .A(grid[320]), .S(n25685), .Y(n27847) );
  MUX2X1 U18226 ( .B(n25605), .A(grid[308]), .S(n27907), .Y(n27851) );
  MUX2X1 U18227 ( .B(n25610), .A(grid[296]), .S(n27910), .Y(n27850) );
  MUX2X1 U18228 ( .B(n27849), .A(n27846), .S(n27915), .Y(n27853) );
  MUX2X1 U18229 ( .B(n25465), .A(grid[284]), .S(n25685), .Y(n27857) );
  MUX2X1 U18230 ( .B(n25598), .A(grid[272]), .S(n25685), .Y(n27856) );
  MUX2X1 U18231 ( .B(grid[254]), .A(n25602), .S(n25685), .Y(n27860) );
  MUX2X1 U18232 ( .B(n25660), .A(grid[248]), .S(n25685), .Y(n27859) );
  MUX2X1 U18233 ( .B(n27858), .A(n27855), .S(n27914), .Y(n27869) );
  MUX2X1 U18234 ( .B(n25509), .A(grid[236]), .S(n25685), .Y(n27863) );
  MUX2X1 U18235 ( .B(grid[218]), .A(grid[224]), .S(n25685), .Y(n27862) );
  MUX2X1 U18236 ( .B(n25654), .A(grid[212]), .S(n25685), .Y(n27866) );
  MUX2X1 U18237 ( .B(n25599), .A(n25499), .S(n25685), .Y(n27865) );
  MUX2X1 U18238 ( .B(n27864), .A(n27861), .S(n27914), .Y(n27868) );
  MUX2X1 U18239 ( .B(n27867), .A(n27852), .S(n25688), .Y(n27901) );
  MUX2X1 U18240 ( .B(grid[182]), .A(grid[188]), .S(n25685), .Y(n27872) );
  MUX2X1 U18241 ( .B(grid[170]), .A(grid[176]), .S(n25685), .Y(n27871) );
  MUX2X1 U18242 ( .B(n25595), .A(grid[164]), .S(n25685), .Y(n27875) );
  MUX2X1 U18243 ( .B(n25574), .A(grid[152]), .S(n25685), .Y(n27874) );
  MUX2X1 U18244 ( .B(n27873), .A(n27870), .S(n27914), .Y(n27884) );
  MUX2X1 U18245 ( .B(grid[134]), .A(grid[140]), .S(n25711), .Y(n27878) );
  MUX2X1 U18246 ( .B(grid[122]), .A(grid[128]), .S(n25711), .Y(n27877) );
  MUX2X1 U18247 ( .B(n25601), .A(grid[116]), .S(n25711), .Y(n27881) );
  MUX2X1 U18248 ( .B(n25495), .A(grid[104]), .S(n25711), .Y(n27880) );
  MUX2X1 U18249 ( .B(n27879), .A(n27876), .S(n27914), .Y(n27883) );
  MUX2X1 U18250 ( .B(grid[86]), .A(grid[92]), .S(n25711), .Y(n27887) );
  MUX2X1 U18251 ( .B(n25503), .A(grid[80]), .S(n25711), .Y(n27886) );
  MUX2X1 U18252 ( .B(n25659), .A(grid[68]), .S(n25711), .Y(n27890) );
  MUX2X1 U18253 ( .B(n25655), .A(n25581), .S(n25711), .Y(n27889) );
  MUX2X1 U18254 ( .B(n27888), .A(n27885), .S(n27914), .Y(n27899) );
  MUX2X1 U18255 ( .B(n25508), .A(grid[44]), .S(n25711), .Y(n27893) );
  MUX2X1 U18256 ( .B(n25484), .A(grid[32]), .S(n25711), .Y(n27892) );
  MUX2X1 U18257 ( .B(n25656), .A(n25582), .S(n25711), .Y(n27896) );
  MUX2X1 U18258 ( .B(n25576), .A(grid[8]), .S(n25711), .Y(n27895) );
  MUX2X1 U18259 ( .B(n27894), .A(n27891), .S(n27914), .Y(n27898) );
  MUX2X1 U18260 ( .B(n27897), .A(n27882), .S(n25619), .Y(n27900) );
  INVX1 U18261 ( .A(n29423), .Y(n27902) );
  MUX2X1 U18262 ( .B(n27919), .A(n27920), .S(net105800), .Y(n27918) );
  MUX2X1 U18263 ( .B(n27922), .A(n27923), .S(net112194), .Y(n27921) );
  MUX2X1 U18264 ( .B(n27925), .A(n27926), .S(net150253), .Y(n27924) );
  MUX2X1 U18265 ( .B(n27928), .A(n27929), .S(net105803), .Y(n27927) );
  MUX2X1 U18266 ( .B(n27931), .A(n27932), .S(n28221), .Y(n27930) );
  MUX2X1 U18267 ( .B(n27934), .A(n27935), .S(net105815), .Y(n27933) );
  MUX2X1 U18268 ( .B(n27937), .A(n27938), .S(net105816), .Y(n27936) );
  MUX2X1 U18269 ( .B(n27940), .A(n27941), .S(net105802), .Y(n27939) );
  MUX2X1 U18270 ( .B(n27943), .A(n27944), .S(net150253), .Y(n27942) );
  MUX2X1 U18271 ( .B(n27946), .A(n27947), .S(n28221), .Y(n27945) );
  MUX2X1 U18272 ( .B(n27949), .A(n27950), .S(net105793), .Y(n27948) );
  MUX2X1 U18273 ( .B(n27952), .A(n27953), .S(net105803), .Y(n27951) );
  MUX2X1 U18274 ( .B(n27955), .A(n27956), .S(net105813), .Y(n27954) );
  MUX2X1 U18275 ( .B(n27958), .A(n27959), .S(net105819), .Y(n27957) );
  MUX2X1 U18276 ( .B(n27961), .A(n27962), .S(n28221), .Y(n27960) );
  MUX2X1 U18277 ( .B(n27964), .A(n27965), .S(net105796), .Y(n27963) );
  MUX2X1 U18278 ( .B(n27967), .A(n27968), .S(net105819), .Y(n27966) );
  MUX2X1 U18279 ( .B(n27970), .A(n27971), .S(net105799), .Y(n27969) );
  MUX2X1 U18280 ( .B(n27973), .A(n27974), .S(net105819), .Y(n27972) );
  MUX2X1 U18281 ( .B(n27976), .A(n27977), .S(n28221), .Y(n27975) );
  MUX2X1 U18282 ( .B(n27979), .A(n27980), .S(net105810), .Y(n27978) );
  MUX2X1 U18283 ( .B(n27982), .A(n27983), .S(net105798), .Y(n27981) );
  MUX2X1 U18284 ( .B(n27985), .A(n27986), .S(net105802), .Y(n27984) );
  MUX2X1 U18285 ( .B(n27988), .A(n27989), .S(net105807), .Y(n27987) );
  MUX2X1 U18286 ( .B(n27994), .A(n27995), .S(net105797), .Y(n27993) );
  MUX2X1 U18287 ( .B(n28000), .A(n28001), .S(net105808), .Y(n27999) );
  MUX2X1 U18288 ( .B(n28003), .A(n28004), .S(net105793), .Y(n28002) );
  MUX2X1 U18289 ( .B(n28006), .A(n28007), .S(n28221), .Y(n28005) );
  MUX2X1 U18290 ( .B(n28009), .A(n28010), .S(net105819), .Y(n28008) );
  MUX2X1 U18291 ( .B(n28012), .A(n28013), .S(net105797), .Y(n28011) );
  MUX2X1 U18292 ( .B(n28018), .A(n28019), .S(net105813), .Y(n28017) );
  MUX2X1 U18293 ( .B(n28024), .A(n28025), .S(net105814), .Y(n28023) );
  MUX2X1 U18294 ( .B(n28027), .A(n28028), .S(net105819), .Y(n28026) );
  MUX2X1 U18295 ( .B(n28041), .A(n28042), .S(net105793), .Y(n28040) );
  MUX2X1 U18296 ( .B(n28047), .A(n28048), .S(net150253), .Y(n28046) );
  MUX2X1 U18297 ( .B(n28056), .A(n28057), .S(net105800), .Y(n28055) );
  MUX2X1 U18298 ( .B(n28065), .A(n28066), .S(net105799), .Y(n28064) );
  MUX2X1 U18299 ( .B(n28068), .A(n28069), .S(n28221), .Y(n28067) );
  MUX2X1 U18300 ( .B(n28071), .A(n28072), .S(net105801), .Y(n28070) );
  MUX2X1 U18301 ( .B(n28074), .A(n28075), .S(net105803), .Y(n28073) );
  MUX2X1 U18302 ( .B(n28077), .A(n28078), .S(net105794), .Y(n28076) );
  MUX2X1 U18303 ( .B(n28086), .A(n28087), .S(net105801), .Y(n28085) );
  MUX2X1 U18304 ( .B(n28089), .A(n28090), .S(net105808), .Y(n28088) );
  MUX2X1 U18305 ( .B(n28092), .A(n28093), .S(net105801), .Y(n28091) );
  MUX2X1 U18306 ( .B(n28098), .A(n28099), .S(n28221), .Y(n28097) );
  MUX2X1 U18307 ( .B(n28101), .A(n28102), .S(net105794), .Y(n28100) );
  MUX2X1 U18308 ( .B(n28104), .A(n28105), .S(net105807), .Y(n28103) );
  MUX2X1 U18309 ( .B(n28107), .A(n28108), .S(net105798), .Y(n28106) );
  MUX2X1 U18310 ( .B(n28110), .A(n28111), .S(net105801), .Y(n28109) );
  MUX2X1 U18311 ( .B(n28113), .A(n28114), .S(net113954), .Y(n28112) );
  MUX2X1 U18312 ( .B(n28116), .A(n28117), .S(net105808), .Y(n28115) );
  MUX2X1 U18313 ( .B(n28119), .A(n28120), .S(net105798), .Y(n28118) );
  MUX2X1 U18314 ( .B(n28122), .A(n28123), .S(net105802), .Y(n28121) );
  MUX2X1 U18315 ( .B(n28125), .A(n28126), .S(net105800), .Y(n28124) );
  MUX2X1 U18316 ( .B(n28131), .A(n28132), .S(net105819), .Y(n28130) );
  MUX2X1 U18317 ( .B(n28134), .A(n28135), .S(net105798), .Y(n28133) );
  MUX2X1 U18318 ( .B(n28137), .A(n28138), .S(net105795), .Y(n28136) );
  MUX2X1 U18319 ( .B(n28140), .A(n28141), .S(net105797), .Y(n28139) );
  MUX2X1 U18320 ( .B(n28143), .A(n28144), .S(n28220), .Y(n28142) );
  MUX2X1 U18321 ( .B(n28146), .A(n28147), .S(net105795), .Y(n28145) );
  MUX2X1 U18322 ( .B(n28149), .A(n28150), .S(net105803), .Y(n28148) );
  MUX2X1 U18323 ( .B(n28152), .A(n28153), .S(net105796), .Y(n28151) );
  MUX2X1 U18324 ( .B(n28155), .A(n28156), .S(net105808), .Y(n28154) );
  MUX2X1 U18325 ( .B(n28158), .A(n28159), .S(n28221), .Y(n28157) );
  MUX2X1 U18326 ( .B(n28173), .A(n28174), .S(net113955), .Y(n28172) );
  MUX2X1 U18327 ( .B(n28176), .A(n28177), .S(net105796), .Y(n28175) );
  MUX2X1 U18328 ( .B(n28182), .A(n28183), .S(net105810), .Y(n28181) );
  MUX2X1 U18329 ( .B(n28185), .A(n28186), .S(net113308), .Y(n28184) );
  MUX2X1 U18330 ( .B(n28188), .A(n28189), .S(net113954), .Y(n28187) );
  MUX2X1 U18331 ( .B(n28191), .A(n28192), .S(net105794), .Y(n28190) );
  MUX2X1 U18332 ( .B(n28194), .A(n28195), .S(net105816), .Y(n28193) );
  MUX2X1 U18333 ( .B(n28197), .A(n28198), .S(net105807), .Y(n28196) );
  MUX2X1 U18334 ( .B(n28203), .A(n28204), .S(net113955), .Y(n28202) );
  MUX2X1 U18335 ( .B(n28206), .A(n28207), .S(net112194), .Y(n28205) );
  MUX2X1 U18336 ( .B(n28209), .A(n28210), .S(net105795), .Y(n28208) );
  MUX2X1 U18337 ( .B(n28212), .A(n28213), .S(net105808), .Y(n28211) );
  MUX2X1 U18338 ( .B(grid[372]), .A(grid[378]), .S(net105859), .Y(n27920) );
  MUX2X1 U18339 ( .B(grid[360]), .A(grid[366]), .S(net116925), .Y(n27919) );
  MUX2X1 U18340 ( .B(grid[348]), .A(grid[354]), .S(alt14_net96238), .Y(n27923)
         );
  MUX2X1 U18341 ( .B(grid[336]), .A(grid[342]), .S(net111222), .Y(n27922) );
  MUX2X1 U18342 ( .B(n27921), .A(n27918), .S(net150046), .Y(n27932) );
  MUX2X1 U18343 ( .B(grid[324]), .A(grid[330]), .S(net151696), .Y(n27926) );
  MUX2X1 U18344 ( .B(grid[312]), .A(grid[318]), .S(net150130), .Y(n27925) );
  MUX2X1 U18345 ( .B(grid[300]), .A(grid[306]), .S(net103671), .Y(n27929) );
  MUX2X1 U18346 ( .B(grid[288]), .A(grid[294]), .S(net151697), .Y(n27928) );
  MUX2X1 U18347 ( .B(n27927), .A(n27924), .S(net149936), .Y(n27931) );
  MUX2X1 U18348 ( .B(grid[276]), .A(grid[282]), .S(net151652), .Y(n27935) );
  MUX2X1 U18349 ( .B(grid[264]), .A(grid[270]), .S(net103671), .Y(n27934) );
  MUX2X1 U18350 ( .B(grid[252]), .A(grid[258]), .S(net103671), .Y(n27938) );
  MUX2X1 U18351 ( .B(grid[240]), .A(grid[246]), .S(net103671), .Y(n27937) );
  MUX2X1 U18352 ( .B(n27936), .A(n27933), .S(net151833), .Y(n27947) );
  MUX2X1 U18353 ( .B(n21088), .A(grid[234]), .S(net147379), .Y(n27941) );
  MUX2X1 U18354 ( .B(grid[216]), .A(grid[222]), .S(net147379), .Y(n27940) );
  MUX2X1 U18355 ( .B(grid[204]), .A(grid[210]), .S(net151652), .Y(n27944) );
  MUX2X1 U18356 ( .B(grid[192]), .A(grid[198]), .S(net105788), .Y(n27943) );
  MUX2X1 U18357 ( .B(n27942), .A(n27939), .S(net149936), .Y(n27946) );
  MUX2X1 U18358 ( .B(grid[180]), .A(grid[186]), .S(net103671), .Y(n27950) );
  MUX2X1 U18359 ( .B(grid[168]), .A(grid[174]), .S(net111222), .Y(n27949) );
  MUX2X1 U18360 ( .B(grid[156]), .A(grid[162]), .S(net150126), .Y(n27953) );
  MUX2X1 U18361 ( .B(grid[144]), .A(grid[150]), .S(net103671), .Y(n27952) );
  MUX2X1 U18362 ( .B(n27951), .A(n27948), .S(net149936), .Y(n27962) );
  MUX2X1 U18363 ( .B(grid[132]), .A(grid[138]), .S(net103671), .Y(n27956) );
  MUX2X1 U18364 ( .B(grid[120]), .A(grid[126]), .S(net103671), .Y(n27955) );
  MUX2X1 U18365 ( .B(grid[108]), .A(grid[114]), .S(net149947), .Y(n27959) );
  MUX2X1 U18366 ( .B(grid[96]), .A(grid[102]), .S(net111222), .Y(n27958) );
  MUX2X1 U18367 ( .B(n27957), .A(n27954), .S(net149936), .Y(n27961) );
  MUX2X1 U18368 ( .B(grid[84]), .A(n21082), .S(net111222), .Y(n27965) );
  MUX2X1 U18369 ( .B(grid[72]), .A(grid[78]), .S(net111222), .Y(n27964) );
  MUX2X1 U18370 ( .B(grid[60]), .A(grid[66]), .S(net103671), .Y(n27968) );
  MUX2X1 U18371 ( .B(grid[48]), .A(grid[54]), .S(net103671), .Y(n27967) );
  MUX2X1 U18372 ( .B(n27966), .A(n27963), .S(net149936), .Y(n27977) );
  MUX2X1 U18373 ( .B(grid[36]), .A(grid[42]), .S(net103671), .Y(n27971) );
  MUX2X1 U18374 ( .B(grid[24]), .A(grid[30]), .S(net105859), .Y(n27970) );
  MUX2X1 U18375 ( .B(grid[12]), .A(grid[18]), .S(net110246), .Y(n27974) );
  MUX2X1 U18376 ( .B(grid[0]), .A(n21086), .S(net103671), .Y(n27973) );
  MUX2X1 U18377 ( .B(n27972), .A(n27969), .S(net149936), .Y(n27976) );
  MUX2X1 U18378 ( .B(grid[373]), .A(grid[379]), .S(net105788), .Y(n27980) );
  MUX2X1 U18379 ( .B(grid[361]), .A(grid[367]), .S(net103671), .Y(n27979) );
  MUX2X1 U18380 ( .B(grid[349]), .A(grid[355]), .S(net114151), .Y(n27983) );
  MUX2X1 U18381 ( .B(grid[337]), .A(grid[343]), .S(net110825), .Y(n27982) );
  MUX2X1 U18382 ( .B(n27981), .A(n27978), .S(net149863), .Y(n27992) );
  MUX2X1 U18383 ( .B(grid[325]), .A(grid[331]), .S(net151697), .Y(n27986) );
  MUX2X1 U18384 ( .B(grid[313]), .A(grid[319]), .S(net105788), .Y(n27985) );
  MUX2X1 U18385 ( .B(grid[301]), .A(grid[307]), .S(net105788), .Y(n27989) );
  MUX2X1 U18386 ( .B(grid[289]), .A(grid[295]), .S(net110246), .Y(n27988) );
  MUX2X1 U18387 ( .B(grid[277]), .A(grid[283]), .S(alt14_net96230), .Y(n27995)
         );
  MUX2X1 U18388 ( .B(grid[265]), .A(grid[271]), .S(net110246), .Y(n27994) );
  MUX2X1 U18389 ( .B(grid[253]), .A(grid[259]), .S(alt14_net96238), .Y(n27998)
         );
  MUX2X1 U18390 ( .B(grid[229]), .A(grid[235]), .S(net110825), .Y(n28001) );
  MUX2X1 U18391 ( .B(grid[217]), .A(grid[223]), .S(net103671), .Y(n28000) );
  MUX2X1 U18392 ( .B(grid[205]), .A(grid[211]), .S(net110825), .Y(n28004) );
  MUX2X1 U18393 ( .B(grid[193]), .A(grid[199]), .S(net110246), .Y(n28003) );
  MUX2X1 U18394 ( .B(n28002), .A(n27999), .S(net149862), .Y(n28006) );
  MUX2X1 U18395 ( .B(n28005), .A(n27990), .S(alt14_net55935), .Y(n28039) );
  MUX2X1 U18396 ( .B(grid[181]), .A(grid[187]), .S(net105788), .Y(n28010) );
  MUX2X1 U18397 ( .B(grid[169]), .A(grid[175]), .S(alt14_net96236), .Y(n28009)
         );
  MUX2X1 U18398 ( .B(n28011), .A(n28008), .S(net151833), .Y(n28022) );
  MUX2X1 U18399 ( .B(grid[121]), .A(grid[127]), .S(net110246), .Y(n28015) );
  MUX2X1 U18400 ( .B(grid[109]), .A(grid[115]), .S(net103671), .Y(n28019) );
  MUX2X1 U18401 ( .B(grid[97]), .A(grid[103]), .S(net116760), .Y(n28018) );
  MUX2X1 U18402 ( .B(n28017), .A(n28014), .S(net149862), .Y(n28021) );
  MUX2X1 U18403 ( .B(grid[85]), .A(grid[91]), .S(net110815), .Y(n28025) );
  MUX2X1 U18404 ( .B(grid[61]), .A(grid[67]), .S(net110815), .Y(n28028) );
  MUX2X1 U18405 ( .B(grid[49]), .A(grid[55]), .S(net105788), .Y(n28027) );
  MUX2X1 U18406 ( .B(n28026), .A(n28023), .S(net149863), .Y(n28037) );
  MUX2X1 U18407 ( .B(grid[25]), .A(grid[31]), .S(net105788), .Y(n28030) );
  MUX2X1 U18408 ( .B(grid[1]), .A(grid[7]), .S(net103671), .Y(n28033) );
  MUX2X1 U18409 ( .B(grid[374]), .A(grid[380]), .S(net111222), .Y(n28042) );
  MUX2X1 U18410 ( .B(grid[362]), .A(grid[368]), .S(alt14_net96230), .Y(n28041)
         );
  MUX2X1 U18411 ( .B(grid[350]), .A(grid[356]), .S(net105788), .Y(n28045) );
  MUX2X1 U18412 ( .B(grid[338]), .A(grid[344]), .S(net111222), .Y(n28044) );
  MUX2X1 U18413 ( .B(n28043), .A(n28040), .S(net149863), .Y(n28054) );
  MUX2X1 U18414 ( .B(grid[326]), .A(grid[332]), .S(net111222), .Y(n28048) );
  MUX2X1 U18415 ( .B(grid[302]), .A(grid[308]), .S(net111222), .Y(n28051) );
  MUX2X1 U18416 ( .B(grid[290]), .A(grid[296]), .S(net110825), .Y(n28050) );
  MUX2X1 U18417 ( .B(n28049), .A(n28046), .S(net149862), .Y(n28053) );
  MUX2X1 U18418 ( .B(grid[278]), .A(grid[284]), .S(net110246), .Y(n28057) );
  MUX2X1 U18419 ( .B(grid[266]), .A(grid[272]), .S(net111222), .Y(n28056) );
  MUX2X1 U18420 ( .B(grid[254]), .A(grid[260]), .S(net114151), .Y(n28060) );
  MUX2X1 U18421 ( .B(n28058), .A(n28055), .S(net151834), .Y(n28069) );
  MUX2X1 U18422 ( .B(grid[218]), .A(grid[224]), .S(net117076), .Y(n28062) );
  MUX2X1 U18423 ( .B(grid[194]), .A(grid[200]), .S(net110246), .Y(n28065) );
  MUX2X1 U18424 ( .B(n28064), .A(n28061), .S(net151833), .Y(n28068) );
  MUX2X1 U18425 ( .B(grid[182]), .A(grid[188]), .S(net103671), .Y(n28072) );
  MUX2X1 U18426 ( .B(grid[170]), .A(grid[176]), .S(net116760), .Y(n28071) );
  MUX2X1 U18427 ( .B(grid[158]), .A(grid[164]), .S(net149947), .Y(n28075) );
  MUX2X1 U18428 ( .B(grid[146]), .A(grid[152]), .S(net151617), .Y(n28074) );
  MUX2X1 U18429 ( .B(n28073), .A(n28070), .S(net151834), .Y(n28084) );
  MUX2X1 U18430 ( .B(grid[134]), .A(grid[140]), .S(net111222), .Y(n28078) );
  MUX2X1 U18431 ( .B(grid[122]), .A(grid[128]), .S(alt14_net96236), .Y(n28077)
         );
  MUX2X1 U18432 ( .B(grid[110]), .A(grid[116]), .S(net149947), .Y(n28081) );
  MUX2X1 U18433 ( .B(grid[98]), .A(grid[104]), .S(net111222), .Y(n28080) );
  MUX2X1 U18434 ( .B(n28079), .A(n28076), .S(net151834), .Y(n28083) );
  MUX2X1 U18435 ( .B(grid[86]), .A(grid[92]), .S(net114151), .Y(n28087) );
  MUX2X1 U18436 ( .B(grid[74]), .A(grid[80]), .S(net114151), .Y(n28086) );
  MUX2X1 U18437 ( .B(grid[50]), .A(grid[56]), .S(net114151), .Y(n28089) );
  MUX2X1 U18438 ( .B(n28088), .A(n28085), .S(net149862), .Y(n28099) );
  MUX2X1 U18439 ( .B(grid[38]), .A(grid[44]), .S(net151696), .Y(n28093) );
  MUX2X1 U18440 ( .B(grid[26]), .A(grid[32]), .S(net116925), .Y(n28092) );
  MUX2X1 U18441 ( .B(grid[14]), .A(grid[20]), .S(net150132), .Y(n28096) );
  MUX2X1 U18442 ( .B(grid[2]), .A(grid[8]), .S(alt14_net96230), .Y(n28095) );
  MUX2X1 U18443 ( .B(n28094), .A(n28091), .S(net151833), .Y(n28098) );
  MUX2X1 U18444 ( .B(n28097), .A(n28082), .S(alt14_net55935), .Y(alt14_net6129) );
  MUX2X1 U18445 ( .B(grid[375]), .A(grid[381]), .S(net105859), .Y(n28102) );
  MUX2X1 U18446 ( .B(grid[363]), .A(grid[369]), .S(net150126), .Y(n28101) );
  MUX2X1 U18447 ( .B(grid[351]), .A(grid[357]), .S(net103671), .Y(n28105) );
  MUX2X1 U18448 ( .B(grid[339]), .A(grid[345]), .S(net111222), .Y(n28104) );
  MUX2X1 U18449 ( .B(n28103), .A(n28100), .S(net149936), .Y(n28114) );
  MUX2X1 U18450 ( .B(grid[327]), .A(grid[333]), .S(net105779), .Y(n28108) );
  MUX2X1 U18451 ( .B(grid[315]), .A(grid[321]), .S(net151617), .Y(n28107) );
  MUX2X1 U18452 ( .B(grid[303]), .A(grid[309]), .S(net147379), .Y(n28111) );
  MUX2X1 U18453 ( .B(grid[291]), .A(grid[297]), .S(net147379), .Y(n28110) );
  MUX2X1 U18454 ( .B(n28109), .A(n28106), .S(net149936), .Y(n28113) );
  MUX2X1 U18455 ( .B(grid[279]), .A(grid[285]), .S(net105859), .Y(n28117) );
  MUX2X1 U18456 ( .B(grid[267]), .A(grid[273]), .S(net150130), .Y(n28116) );
  MUX2X1 U18457 ( .B(grid[255]), .A(grid[261]), .S(net105859), .Y(n28120) );
  MUX2X1 U18458 ( .B(grid[243]), .A(grid[249]), .S(net147379), .Y(n28119) );
  MUX2X1 U18459 ( .B(n28118), .A(n28115), .S(net149936), .Y(n28129) );
  MUX2X1 U18460 ( .B(grid[231]), .A(grid[237]), .S(net105859), .Y(n28123) );
  MUX2X1 U18461 ( .B(grid[207]), .A(grid[213]), .S(net105859), .Y(n28126) );
  MUX2X1 U18462 ( .B(grid[195]), .A(grid[201]), .S(net111222), .Y(n28125) );
  MUX2X1 U18463 ( .B(n28124), .A(n28121), .S(net149936), .Y(n28128) );
  MUX2X1 U18464 ( .B(n28127), .A(n28112), .S(alt14_net55927), .Y(alt14_net6192) );
  MUX2X1 U18465 ( .B(grid[183]), .A(grid[189]), .S(net105859), .Y(n28132) );
  MUX2X1 U18466 ( .B(grid[171]), .A(grid[177]), .S(net105859), .Y(n28131) );
  MUX2X1 U18467 ( .B(grid[159]), .A(grid[165]), .S(net105859), .Y(n28135) );
  MUX2X1 U18468 ( .B(grid[147]), .A(grid[153]), .S(net105859), .Y(n28134) );
  MUX2X1 U18469 ( .B(n28133), .A(n28130), .S(net149936), .Y(n28144) );
  MUX2X1 U18470 ( .B(grid[135]), .A(grid[141]), .S(net105859), .Y(n28138) );
  MUX2X1 U18471 ( .B(grid[123]), .A(grid[129]), .S(net151617), .Y(n28137) );
  MUX2X1 U18472 ( .B(grid[111]), .A(grid[117]), .S(net105859), .Y(n28141) );
  MUX2X1 U18473 ( .B(grid[99]), .A(grid[105]), .S(net105859), .Y(n28140) );
  MUX2X1 U18474 ( .B(n28139), .A(n28136), .S(net149936), .Y(n28143) );
  MUX2X1 U18475 ( .B(grid[87]), .A(grid[93]), .S(net105779), .Y(n28147) );
  MUX2X1 U18476 ( .B(grid[75]), .A(grid[81]), .S(net105779), .Y(n28146) );
  MUX2X1 U18477 ( .B(grid[63]), .A(grid[69]), .S(net105779), .Y(n28150) );
  MUX2X1 U18478 ( .B(grid[51]), .A(grid[57]), .S(net105779), .Y(n28149) );
  MUX2X1 U18479 ( .B(n28148), .A(n28145), .S(net150046), .Y(n28159) );
  MUX2X1 U18480 ( .B(grid[39]), .A(grid[45]), .S(net105779), .Y(n28153) );
  MUX2X1 U18481 ( .B(grid[27]), .A(grid[33]), .S(net105779), .Y(n28152) );
  MUX2X1 U18482 ( .B(grid[15]), .A(grid[21]), .S(net105779), .Y(n28156) );
  MUX2X1 U18483 ( .B(grid[3]), .A(grid[9]), .S(net105779), .Y(n28155) );
  MUX2X1 U18484 ( .B(n28154), .A(n28151), .S(net149863), .Y(n28158) );
  MUX2X1 U18485 ( .B(n28157), .A(n28142), .S(alt14_net55927), .Y(alt14_net6191) );
  MUX2X1 U18486 ( .B(grid[340]), .A(grid[346]), .S(net112202), .Y(n28164) );
  MUX2X1 U18487 ( .B(grid[316]), .A(grid[322]), .S(alt14_net96236), .Y(n28167)
         );
  MUX2X1 U18488 ( .B(grid[292]), .A(grid[298]), .S(alt14_net96236), .Y(n28170)
         );
  MUX2X1 U18489 ( .B(n28169), .A(n28166), .S(net149936), .Y(n28173) );
  MUX2X1 U18490 ( .B(grid[280]), .A(grid[286]), .S(alt14_net96236), .Y(n28177)
         );
  MUX2X1 U18491 ( .B(grid[268]), .A(grid[274]), .S(n20807), .Y(n28176) );
  MUX2X1 U18492 ( .B(grid[244]), .A(grid[250]), .S(net110825), .Y(n28179) );
  MUX2X1 U18493 ( .B(grid[232]), .A(grid[238]), .S(net105788), .Y(n28183) );
  MUX2X1 U18494 ( .B(grid[208]), .A(grid[214]), .S(net112202), .Y(n28186) );
  MUX2X1 U18495 ( .B(grid[196]), .A(grid[202]), .S(net112202), .Y(n28185) );
  MUX2X1 U18496 ( .B(n28184), .A(n28181), .S(net149936), .Y(n28188) );
  MUX2X1 U18497 ( .B(grid[184]), .A(grid[190]), .S(net105788), .Y(n28192) );
  MUX2X1 U18498 ( .B(grid[172]), .A(grid[178]), .S(net110246), .Y(n28191) );
  MUX2X1 U18499 ( .B(grid[160]), .A(grid[166]), .S(net112202), .Y(n28195) );
  MUX2X1 U18500 ( .B(grid[148]), .A(grid[154]), .S(net112202), .Y(n28194) );
  MUX2X1 U18501 ( .B(n28193), .A(n28190), .S(net149986), .Y(n28204) );
  MUX2X1 U18502 ( .B(grid[136]), .A(grid[142]), .S(alt14_net96236), .Y(n28198)
         );
  MUX2X1 U18503 ( .B(grid[124]), .A(grid[130]), .S(net110246), .Y(n28197) );
  MUX2X1 U18504 ( .B(grid[112]), .A(grid[118]), .S(alt14_net96236), .Y(n28201)
         );
  MUX2X1 U18505 ( .B(grid[100]), .A(grid[106]), .S(alt14_net96236), .Y(n28200)
         );
  MUX2X1 U18506 ( .B(n28199), .A(n28196), .S(net149986), .Y(n28203) );
  MUX2X1 U18507 ( .B(grid[88]), .A(grid[94]), .S(alt14_net96230), .Y(n28207)
         );
  MUX2X1 U18508 ( .B(grid[52]), .A(grid[58]), .S(alt14_net96230), .Y(n28209)
         );
  MUX2X1 U18509 ( .B(n28208), .A(n28205), .S(net149986), .Y(n28219) );
  MUX2X1 U18510 ( .B(grid[40]), .A(grid[46]), .S(net112202), .Y(n28213) );
  MUX2X1 U18511 ( .B(grid[28]), .A(grid[34]), .S(net112202), .Y(n28212) );
  MUX2X1 U18512 ( .B(grid[4]), .A(grid[10]), .S(net105787), .Y(n28215) );
  MUX2X1 U18513 ( .B(n28214), .A(n28211), .S(net149986), .Y(n28218) );
  MUX2X1 U18514 ( .B(n28217), .A(n28202), .S(alt14_net55921), .Y(alt14_net6253) );
  MUX2X1 U18515 ( .B(n28223), .A(n28224), .S(n26486), .Y(n28222) );
  MUX2X1 U18516 ( .B(n28226), .A(n28227), .S(n26513), .Y(n28225) );
  MUX2X1 U18517 ( .B(n28229), .A(n28230), .S(n26505), .Y(n28228) );
  MUX2X1 U18518 ( .B(n28232), .A(n28233), .S(n26505), .Y(n28231) );
  MUX2X1 U18519 ( .B(n28235), .A(n28236), .S(n28607), .Y(n28234) );
  MUX2X1 U18520 ( .B(n28238), .A(n28239), .S(n26512), .Y(n28237) );
  MUX2X1 U18521 ( .B(n28241), .A(n28242), .S(n26503), .Y(n28240) );
  MUX2X1 U18522 ( .B(n28244), .A(n28245), .S(n26506), .Y(n28243) );
  MUX2X1 U18523 ( .B(n28247), .A(n28248), .S(n26509), .Y(n28246) );
  MUX2X1 U18524 ( .B(n28250), .A(n28251), .S(n28607), .Y(n28249) );
  MUX2X1 U18525 ( .B(n28253), .A(n28254), .S(n26488), .Y(n28252) );
  MUX2X1 U18526 ( .B(n28256), .A(n28257), .S(n26487), .Y(n28255) );
  MUX2X1 U18527 ( .B(n28262), .A(n28263), .S(n26486), .Y(n28261) );
  MUX2X1 U18528 ( .B(n28265), .A(n28266), .S(n28607), .Y(n28264) );
  MUX2X1 U18529 ( .B(n28268), .A(n28269), .S(n26490), .Y(n28267) );
  MUX2X1 U18530 ( .B(n28271), .A(n28272), .S(n26492), .Y(n28270) );
  MUX2X1 U18531 ( .B(n28274), .A(n28275), .S(n26486), .Y(n28273) );
  MUX2X1 U18532 ( .B(n28277), .A(n28278), .S(n26486), .Y(n28276) );
  MUX2X1 U18533 ( .B(n28280), .A(n28281), .S(n28607), .Y(n28279) );
  MUX2X1 U18534 ( .B(n28282), .A(n28283), .S(n27211), .Y(n8039) );
  MUX2X1 U18535 ( .B(n28285), .A(n28286), .S(n26511), .Y(n28284) );
  MUX2X1 U18536 ( .B(n28288), .A(n28289), .S(n26499), .Y(n28287) );
  MUX2X1 U18537 ( .B(n28291), .A(n28292), .S(n26511), .Y(n28290) );
  MUX2X1 U18538 ( .B(n28294), .A(n28295), .S(n26492), .Y(n28293) );
  MUX2X1 U18539 ( .B(n28297), .A(n28298), .S(n28607), .Y(n28296) );
  MUX2X1 U18540 ( .B(n28300), .A(n28301), .S(n26498), .Y(n28299) );
  MUX2X1 U18541 ( .B(n28303), .A(n28304), .S(n26501), .Y(n28302) );
  MUX2X1 U18542 ( .B(n28306), .A(n28307), .S(n26500), .Y(n28305) );
  MUX2X1 U18543 ( .B(n28309), .A(n28310), .S(n26489), .Y(n28308) );
  MUX2X1 U18544 ( .B(n28312), .A(n28313), .S(n28607), .Y(n28311) );
  MUX2X1 U18545 ( .B(n28315), .A(n28316), .S(n26510), .Y(n28314) );
  MUX2X1 U18546 ( .B(n28318), .A(n28319), .S(n26508), .Y(n28317) );
  MUX2X1 U18547 ( .B(n28324), .A(n28325), .S(n26486), .Y(n28323) );
  MUX2X1 U18548 ( .B(n28330), .A(n28331), .S(n26508), .Y(n28329) );
  MUX2X1 U18549 ( .B(n28333), .A(n28334), .S(n26500), .Y(n28332) );
  MUX2X1 U18550 ( .B(n28336), .A(n28337), .S(n26495), .Y(n28335) );
  MUX2X1 U18551 ( .B(n28339), .A(n28340), .S(n26494), .Y(n28338) );
  MUX2X1 U18552 ( .B(n28342), .A(n28343), .S(n28607), .Y(n28341) );
  MUX2X1 U18553 ( .B(n28344), .A(n28345), .S(n27210), .Y(n8038) );
  MUX2X1 U18554 ( .B(n28347), .A(n28348), .S(n26501), .Y(n28346) );
  MUX2X1 U18555 ( .B(n28350), .A(n28351), .S(n26506), .Y(n28349) );
  MUX2X1 U18556 ( .B(n28353), .A(n28354), .S(n26493), .Y(n28352) );
  MUX2X1 U18557 ( .B(n28356), .A(n28357), .S(n26486), .Y(n28355) );
  MUX2X1 U18558 ( .B(n28359), .A(n28360), .S(n28607), .Y(n28358) );
  MUX2X1 U18559 ( .B(n28362), .A(n28363), .S(n26504), .Y(n28361) );
  MUX2X1 U18560 ( .B(n28368), .A(n28369), .S(n26513), .Y(n28367) );
  MUX2X1 U18561 ( .B(n28371), .A(n28372), .S(n26490), .Y(n28370) );
  MUX2X1 U18562 ( .B(n28374), .A(n28375), .S(n28607), .Y(n28373) );
  MUX2X1 U18563 ( .B(n28377), .A(n28378), .S(n26504), .Y(n28376) );
  MUX2X1 U18564 ( .B(n28380), .A(n28381), .S(n26512), .Y(n28379) );
  MUX2X1 U18565 ( .B(n28383), .A(n28384), .S(n26498), .Y(n28382) );
  MUX2X1 U18566 ( .B(n28386), .A(n28387), .S(n26495), .Y(n28385) );
  MUX2X1 U18567 ( .B(n28389), .A(n28390), .S(n28607), .Y(n28388) );
  MUX2X1 U18568 ( .B(n28392), .A(n28393), .S(n21043), .Y(n28391) );
  MUX2X1 U18569 ( .B(n28395), .A(n28396), .S(n26489), .Y(n28394) );
  MUX2X1 U18570 ( .B(n28398), .A(n28399), .S(n26494), .Y(n28397) );
  MUX2X1 U18571 ( .B(n28401), .A(n28402), .S(n26487), .Y(n28400) );
  MUX2X1 U18572 ( .B(n28404), .A(n28405), .S(n28607), .Y(n28403) );
  MUX2X1 U18573 ( .B(n28406), .A(n28407), .S(n27210), .Y(n8037) );
  MUX2X1 U18574 ( .B(n28409), .A(n28410), .S(n26502), .Y(n28408) );
  MUX2X1 U18575 ( .B(n28412), .A(n28413), .S(n26488), .Y(n28411) );
  MUX2X1 U18576 ( .B(n28415), .A(n28416), .S(n26497), .Y(n28414) );
  MUX2X1 U18577 ( .B(n28418), .A(n28419), .S(n26490), .Y(n28417) );
  MUX2X1 U18578 ( .B(n28421), .A(n28422), .S(n28606), .Y(n28420) );
  MUX2X1 U18579 ( .B(n28424), .A(n28425), .S(n26491), .Y(n28423) );
  MUX2X1 U18580 ( .B(n28427), .A(n28428), .S(n26507), .Y(n28426) );
  MUX2X1 U18581 ( .B(n28430), .A(n28431), .S(n26489), .Y(n28429) );
  MUX2X1 U18582 ( .B(n28433), .A(n28434), .S(n26492), .Y(n28432) );
  MUX2X1 U18583 ( .B(n28436), .A(n28437), .S(n28606), .Y(n28435) );
  MUX2X1 U18584 ( .B(n28439), .A(n28440), .S(n26496), .Y(n28438) );
  MUX2X1 U18585 ( .B(n28442), .A(n28443), .S(n26488), .Y(n28441) );
  MUX2X1 U18586 ( .B(n28445), .A(n28446), .S(n26487), .Y(n28444) );
  MUX2X1 U18587 ( .B(n28448), .A(n28449), .S(n26500), .Y(n28447) );
  MUX2X1 U18588 ( .B(n28451), .A(n28452), .S(n28606), .Y(n28450) );
  MUX2X1 U18589 ( .B(n28454), .A(n28455), .S(n26487), .Y(n28453) );
  MUX2X1 U18590 ( .B(n28460), .A(n28461), .S(n26499), .Y(n28459) );
  MUX2X1 U18591 ( .B(n28463), .A(n28464), .S(n26504), .Y(n28462) );
  MUX2X1 U18592 ( .B(n28466), .A(n28467), .S(n28606), .Y(n28465) );
  MUX2X1 U18593 ( .B(n28468), .A(n28469), .S(n27210), .Y(n8036) );
  MUX2X1 U18594 ( .B(n28471), .A(n28472), .S(n26503), .Y(n28470) );
  MUX2X1 U18595 ( .B(n28477), .A(n28478), .S(n26489), .Y(n28476) );
  MUX2X1 U18596 ( .B(n28483), .A(n28484), .S(n28606), .Y(n28482) );
  MUX2X1 U18597 ( .B(n28489), .A(n28490), .S(n26491), .Y(n28488) );
  MUX2X1 U18598 ( .B(n28495), .A(n28496), .S(n26493), .Y(n28494) );
  MUX2X1 U18599 ( .B(n28498), .A(n28499), .S(n28607), .Y(n28497) );
  MUX2X1 U18600 ( .B(n28501), .A(n28502), .S(n26497), .Y(n28500) );
  MUX2X1 U18601 ( .B(n28504), .A(n28505), .S(n26490), .Y(n28503) );
  MUX2X1 U18602 ( .B(n28510), .A(n28511), .S(n26496), .Y(n28509) );
  MUX2X1 U18603 ( .B(n28516), .A(n28517), .S(n26489), .Y(n28515) );
  MUX2X1 U18604 ( .B(n28519), .A(n28520), .S(n26494), .Y(n28518) );
  MUX2X1 U18605 ( .B(n28522), .A(n28523), .S(n26495), .Y(n28521) );
  MUX2X1 U18606 ( .B(n28528), .A(n28529), .S(n28606), .Y(n28527) );
  MUX2X1 U18607 ( .B(n28530), .A(n28531), .S(n27209), .Y(n8035) );
  MUX2X1 U18608 ( .B(n28533), .A(n28534), .S(n26510), .Y(n28532) );
  MUX2X1 U18609 ( .B(n28536), .A(n28537), .S(n26488), .Y(n28535) );
  MUX2X1 U18610 ( .B(n28539), .A(n28540), .S(n26498), .Y(n28538) );
  MUX2X1 U18611 ( .B(n28542), .A(n28543), .S(n26502), .Y(n28541) );
  MUX2X1 U18612 ( .B(n28545), .A(n28546), .S(n28606), .Y(n28544) );
  MUX2X1 U18613 ( .B(n28548), .A(n28549), .S(n26487), .Y(n28547) );
  MUX2X1 U18614 ( .B(n28551), .A(n28552), .S(n26488), .Y(n28550) );
  MUX2X1 U18615 ( .B(n28554), .A(n28555), .S(n26490), .Y(n28553) );
  MUX2X1 U18616 ( .B(n28557), .A(n28558), .S(n26496), .Y(n28556) );
  MUX2X1 U18617 ( .B(n28563), .A(n28564), .S(n26499), .Y(n28562) );
  MUX2X1 U18618 ( .B(n28566), .A(n28567), .S(n21043), .Y(n28565) );
  MUX2X1 U18619 ( .B(n28569), .A(n28570), .S(n26492), .Y(n28568) );
  MUX2X1 U18620 ( .B(n28572), .A(n28573), .S(n26492), .Y(n28571) );
  MUX2X1 U18621 ( .B(n28575), .A(n28576), .S(n28606), .Y(n28574) );
  MUX2X1 U18622 ( .B(n28578), .A(n28579), .S(n26504), .Y(n28577) );
  MUX2X1 U18623 ( .B(n28581), .A(n28582), .S(n26506), .Y(n28580) );
  MUX2X1 U18624 ( .B(n28587), .A(n28588), .S(n26493), .Y(n28586) );
  MUX2X1 U18625 ( .B(n28590), .A(n28591), .S(n28606), .Y(n28589) );
  MUX2X1 U18626 ( .B(n28592), .A(n28593), .S(n27209), .Y(n8034) );
  MUX2X1 U18627 ( .B(grid[372]), .A(grid[378]), .S(n26123), .Y(n28224) );
  MUX2X1 U18628 ( .B(grid[360]), .A(grid[366]), .S(n26136), .Y(n28223) );
  MUX2X1 U18629 ( .B(n25626), .A(grid[354]), .S(n26124), .Y(n28227) );
  MUX2X1 U18630 ( .B(grid[336]), .A(grid[342]), .S(n26130), .Y(n28226) );
  MUX2X1 U18631 ( .B(n28225), .A(n28222), .S(n29462), .Y(n28236) );
  MUX2X1 U18632 ( .B(grid[324]), .A(grid[330]), .S(n26081), .Y(n28230) );
  MUX2X1 U18633 ( .B(grid[312]), .A(grid[318]), .S(n26109), .Y(n28229) );
  MUX2X1 U18634 ( .B(n25618), .A(grid[306]), .S(n26138), .Y(n28233) );
  MUX2X1 U18635 ( .B(grid[288]), .A(grid[294]), .S(n26121), .Y(n28232) );
  MUX2X1 U18636 ( .B(n28231), .A(n28228), .S(n29462), .Y(n28235) );
  MUX2X1 U18637 ( .B(grid[276]), .A(grid[282]), .S(n26125), .Y(n28239) );
  MUX2X1 U18638 ( .B(grid[264]), .A(grid[270]), .S(n26083), .Y(n28238) );
  MUX2X1 U18639 ( .B(n25643), .A(grid[258]), .S(n26126), .Y(n28242) );
  MUX2X1 U18640 ( .B(n25637), .A(grid[246]), .S(n26148), .Y(n28241) );
  MUX2X1 U18641 ( .B(n21088), .A(grid[234]), .S(n26138), .Y(n28245) );
  MUX2X1 U18642 ( .B(grid[216]), .A(grid[222]), .S(n26084), .Y(n28244) );
  MUX2X1 U18643 ( .B(n25635), .A(grid[210]), .S(n26089), .Y(n28248) );
  MUX2X1 U18644 ( .B(n25631), .A(grid[198]), .S(n26104), .Y(n28247) );
  MUX2X1 U18645 ( .B(n28246), .A(n28243), .S(n29462), .Y(n28250) );
  MUX2X1 U18646 ( .B(n28249), .A(n28234), .S(n28608), .Y(n28283) );
  MUX2X1 U18647 ( .B(grid[180]), .A(grid[186]), .S(n26079), .Y(n28254) );
  MUX2X1 U18648 ( .B(grid[168]), .A(grid[174]), .S(n26133), .Y(n28253) );
  MUX2X1 U18649 ( .B(grid[156]), .A(grid[162]), .S(n26137), .Y(n28257) );
  MUX2X1 U18650 ( .B(n21084), .A(grid[150]), .S(n26086), .Y(n28256) );
  MUX2X1 U18651 ( .B(n28255), .A(n28252), .S(n26304), .Y(n28266) );
  MUX2X1 U18652 ( .B(grid[132]), .A(grid[138]), .S(n26118), .Y(n28260) );
  MUX2X1 U18653 ( .B(grid[120]), .A(grid[126]), .S(n26088), .Y(n28259) );
  MUX2X1 U18654 ( .B(grid[108]), .A(grid[114]), .S(n26091), .Y(n28263) );
  MUX2X1 U18655 ( .B(grid[96]), .A(grid[102]), .S(n26091), .Y(n28262) );
  MUX2X1 U18656 ( .B(n28261), .A(n28258), .S(n29462), .Y(n28265) );
  MUX2X1 U18657 ( .B(grid[84]), .A(n21082), .S(n26086), .Y(n28269) );
  MUX2X1 U18658 ( .B(grid[72]), .A(grid[78]), .S(n26119), .Y(n28268) );
  MUX2X1 U18659 ( .B(n25639), .A(grid[66]), .S(n26091), .Y(n28272) );
  MUX2X1 U18660 ( .B(grid[48]), .A(grid[54]), .S(n26117), .Y(n28271) );
  MUX2X1 U18661 ( .B(n28270), .A(n28267), .S(n29462), .Y(n28281) );
  MUX2X1 U18662 ( .B(grid[36]), .A(grid[42]), .S(n26092), .Y(n28275) );
  MUX2X1 U18663 ( .B(grid[24]), .A(grid[30]), .S(n26119), .Y(n28274) );
  MUX2X1 U18664 ( .B(grid[12]), .A(grid[18]), .S(n26100), .Y(n28278) );
  MUX2X1 U18665 ( .B(grid[0]), .A(n21086), .S(n26092), .Y(n28277) );
  MUX2X1 U18666 ( .B(n28276), .A(n28273), .S(n26304), .Y(n28280) );
  MUX2X1 U18667 ( .B(n28279), .A(n28264), .S(n28608), .Y(n28282) );
  MUX2X1 U18668 ( .B(grid[373]), .A(grid[379]), .S(n26105), .Y(n28286) );
  MUX2X1 U18669 ( .B(grid[361]), .A(n21215), .S(n26136), .Y(n28285) );
  MUX2X1 U18670 ( .B(grid[349]), .A(grid[355]), .S(n26094), .Y(n28289) );
  MUX2X1 U18671 ( .B(grid[337]), .A(grid[343]), .S(n26132), .Y(n28288) );
  MUX2X1 U18672 ( .B(n28287), .A(n28284), .S(n26304), .Y(n28298) );
  MUX2X1 U18673 ( .B(grid[325]), .A(n23205), .S(n26141), .Y(n28292) );
  MUX2X1 U18674 ( .B(grid[313]), .A(grid[319]), .S(n20847), .Y(n28291) );
  MUX2X1 U18675 ( .B(grid[301]), .A(n25493), .S(n26114), .Y(n28295) );
  MUX2X1 U18676 ( .B(grid[289]), .A(grid[295]), .S(n26106), .Y(n28294) );
  MUX2X1 U18677 ( .B(n28293), .A(n28290), .S(n29462), .Y(n28297) );
  MUX2X1 U18678 ( .B(n25513), .A(grid[283]), .S(n26108), .Y(n28301) );
  MUX2X1 U18679 ( .B(n25506), .A(grid[271]), .S(n26090), .Y(n28300) );
  MUX2X1 U18680 ( .B(grid[253]), .A(grid[259]), .S(n26082), .Y(n28304) );
  MUX2X1 U18681 ( .B(n25487), .A(n25494), .S(n26127), .Y(n28303) );
  MUX2X1 U18682 ( .B(n28302), .A(n28299), .S(n29462), .Y(n28313) );
  MUX2X1 U18683 ( .B(grid[229]), .A(grid[235]), .S(n26131), .Y(n28307) );
  MUX2X1 U18684 ( .B(grid[217]), .A(n20831), .S(n26099), .Y(n28306) );
  MUX2X1 U18685 ( .B(n25600), .A(grid[211]), .S(n26126), .Y(n28310) );
  MUX2X1 U18686 ( .B(grid[193]), .A(grid[199]), .S(n26147), .Y(n28309) );
  MUX2X1 U18687 ( .B(n28308), .A(n28305), .S(n26304), .Y(n28312) );
  MUX2X1 U18688 ( .B(n28311), .A(n28296), .S(n28608), .Y(n28345) );
  MUX2X1 U18689 ( .B(grid[181]), .A(n25496), .S(n26129), .Y(n28316) );
  MUX2X1 U18690 ( .B(grid[169]), .A(grid[175]), .S(n26104), .Y(n28315) );
  MUX2X1 U18691 ( .B(grid[157]), .A(grid[163]), .S(n26087), .Y(n28319) );
  MUX2X1 U18692 ( .B(grid[145]), .A(grid[151]), .S(n26110), .Y(n28318) );
  MUX2X1 U18693 ( .B(n28317), .A(n28314), .S(n29462), .Y(n28328) );
  MUX2X1 U18694 ( .B(grid[133]), .A(grid[139]), .S(n26116), .Y(n28322) );
  MUX2X1 U18695 ( .B(grid[121]), .A(grid[127]), .S(n26096), .Y(n28321) );
  MUX2X1 U18696 ( .B(grid[109]), .A(grid[115]), .S(n26098), .Y(n28325) );
  MUX2X1 U18697 ( .B(n28323), .A(n28320), .S(n26304), .Y(n28327) );
  MUX2X1 U18698 ( .B(grid[85]), .A(n25501), .S(n26148), .Y(n28331) );
  MUX2X1 U18699 ( .B(n25578), .A(grid[79]), .S(n26100), .Y(n28330) );
  MUX2X1 U18700 ( .B(grid[61]), .A(grid[67]), .S(n26113), .Y(n28334) );
  MUX2X1 U18701 ( .B(grid[49]), .A(grid[55]), .S(n26146), .Y(n28333) );
  MUX2X1 U18702 ( .B(n28332), .A(n28329), .S(n29462), .Y(n28343) );
  MUX2X1 U18703 ( .B(n25511), .A(grid[43]), .S(n26097), .Y(n28337) );
  MUX2X1 U18704 ( .B(grid[13]), .A(grid[19]), .S(n26145), .Y(n28340) );
  MUX2X1 U18705 ( .B(grid[1]), .A(grid[7]), .S(n26133), .Y(n28339) );
  MUX2X1 U18706 ( .B(n28338), .A(n28335), .S(n29462), .Y(n28342) );
  MUX2X1 U18707 ( .B(grid[374]), .A(grid[380]), .S(n26161), .Y(n28348) );
  MUX2X1 U18708 ( .B(grid[362]), .A(grid[368]), .S(n26092), .Y(n28347) );
  MUX2X1 U18709 ( .B(grid[350]), .A(grid[356]), .S(n26102), .Y(n28351) );
  MUX2X1 U18710 ( .B(n25500), .A(grid[344]), .S(n26082), .Y(n28350) );
  MUX2X1 U18711 ( .B(n28349), .A(n28346), .S(n26304), .Y(n28360) );
  MUX2X1 U18712 ( .B(n25502), .A(grid[332]), .S(n26096), .Y(n28354) );
  MUX2X1 U18713 ( .B(grid[314]), .A(grid[320]), .S(n26110), .Y(n28353) );
  MUX2X1 U18714 ( .B(n25605), .A(grid[308]), .S(n26083), .Y(n28357) );
  MUX2X1 U18715 ( .B(n25610), .A(grid[296]), .S(n26115), .Y(n28356) );
  MUX2X1 U18716 ( .B(n28355), .A(n28352), .S(n29462), .Y(n28359) );
  MUX2X1 U18717 ( .B(n25465), .A(grid[284]), .S(n26116), .Y(n28363) );
  MUX2X1 U18718 ( .B(n25598), .A(grid[272]), .S(n26085), .Y(n28362) );
  MUX2X1 U18719 ( .B(grid[254]), .A(n25602), .S(n26127), .Y(n28366) );
  MUX2X1 U18720 ( .B(n25660), .A(grid[248]), .S(n26158), .Y(n28365) );
  MUX2X1 U18721 ( .B(n28364), .A(n28361), .S(n26304), .Y(n28375) );
  MUX2X1 U18722 ( .B(n25509), .A(grid[236]), .S(n26155), .Y(n28369) );
  MUX2X1 U18723 ( .B(grid[218]), .A(grid[224]), .S(n26107), .Y(n28368) );
  MUX2X1 U18724 ( .B(grid[206]), .A(grid[212]), .S(n26159), .Y(n28372) );
  MUX2X1 U18725 ( .B(n25505), .A(grid[200]), .S(n26120), .Y(n28371) );
  MUX2X1 U18726 ( .B(n28370), .A(n28367), .S(n29462), .Y(n28374) );
  MUX2X1 U18727 ( .B(n28373), .A(n28358), .S(n28608), .Y(n28407) );
  MUX2X1 U18728 ( .B(grid[182]), .A(grid[188]), .S(n26081), .Y(n28378) );
  MUX2X1 U18729 ( .B(grid[170]), .A(grid[176]), .S(n26098), .Y(n28377) );
  MUX2X1 U18730 ( .B(n25595), .A(grid[164]), .S(n26087), .Y(n28381) );
  MUX2X1 U18731 ( .B(n25574), .A(grid[152]), .S(n26116), .Y(n28380) );
  MUX2X1 U18732 ( .B(n28379), .A(n28376), .S(n21129), .Y(n28390) );
  MUX2X1 U18733 ( .B(grid[134]), .A(grid[140]), .S(n26099), .Y(n28384) );
  MUX2X1 U18734 ( .B(grid[122]), .A(grid[128]), .S(n26127), .Y(n28383) );
  MUX2X1 U18735 ( .B(n25601), .A(grid[116]), .S(n26118), .Y(n28387) );
  MUX2X1 U18736 ( .B(n25495), .A(grid[104]), .S(n26080), .Y(n28386) );
  MUX2X1 U18737 ( .B(n28385), .A(n28382), .S(n29462), .Y(n28389) );
  MUX2X1 U18738 ( .B(grid[86]), .A(grid[92]), .S(n26154), .Y(n28393) );
  MUX2X1 U18739 ( .B(n25503), .A(grid[80]), .S(n26108), .Y(n28392) );
  MUX2X1 U18740 ( .B(n25659), .A(grid[68]), .S(n26160), .Y(n28396) );
  MUX2X1 U18741 ( .B(n25655), .A(grid[56]), .S(n26087), .Y(n28395) );
  MUX2X1 U18742 ( .B(n28394), .A(n28391), .S(n29462), .Y(n28405) );
  MUX2X1 U18743 ( .B(n25508), .A(grid[44]), .S(n26135), .Y(n28399) );
  MUX2X1 U18744 ( .B(n25484), .A(grid[32]), .S(n26080), .Y(n28398) );
  MUX2X1 U18745 ( .B(n25656), .A(grid[20]), .S(n26114), .Y(n28402) );
  MUX2X1 U18746 ( .B(n25576), .A(grid[8]), .S(n26102), .Y(n28401) );
  MUX2X1 U18747 ( .B(n28400), .A(n28397), .S(n29462), .Y(n28404) );
  MUX2X1 U18748 ( .B(grid[375]), .A(grid[381]), .S(n26109), .Y(n28410) );
  MUX2X1 U18749 ( .B(grid[363]), .A(grid[369]), .S(n26134), .Y(n28409) );
  MUX2X1 U18750 ( .B(grid[351]), .A(grid[357]), .S(n26140), .Y(n28413) );
  MUX2X1 U18751 ( .B(grid[339]), .A(grid[345]), .S(n26156), .Y(n28412) );
  MUX2X1 U18752 ( .B(n28411), .A(n28408), .S(n29462), .Y(n28422) );
  MUX2X1 U18753 ( .B(grid[327]), .A(grid[333]), .S(n26152), .Y(n28416) );
  MUX2X1 U18754 ( .B(grid[315]), .A(grid[321]), .S(n26111), .Y(n28415) );
  MUX2X1 U18755 ( .B(grid[303]), .A(grid[309]), .S(n26157), .Y(n28419) );
  MUX2X1 U18756 ( .B(grid[291]), .A(grid[297]), .S(n26090), .Y(n28418) );
  MUX2X1 U18757 ( .B(n28417), .A(n28414), .S(n29462), .Y(n28421) );
  MUX2X1 U18758 ( .B(grid[279]), .A(grid[285]), .S(n26084), .Y(n28425) );
  MUX2X1 U18759 ( .B(grid[267]), .A(grid[273]), .S(n26105), .Y(n28424) );
  MUX2X1 U18760 ( .B(grid[255]), .A(grid[261]), .S(n26122), .Y(n28428) );
  MUX2X1 U18761 ( .B(grid[243]), .A(grid[249]), .S(n26117), .Y(n28427) );
  MUX2X1 U18762 ( .B(n28426), .A(n28423), .S(n26304), .Y(n28437) );
  MUX2X1 U18763 ( .B(grid[231]), .A(grid[237]), .S(n26154), .Y(n28431) );
  MUX2X1 U18764 ( .B(grid[219]), .A(grid[225]), .S(n26084), .Y(n28430) );
  MUX2X1 U18765 ( .B(grid[207]), .A(grid[213]), .S(n26115), .Y(n28434) );
  MUX2X1 U18766 ( .B(grid[195]), .A(grid[201]), .S(n26130), .Y(n28433) );
  MUX2X1 U18767 ( .B(n28432), .A(n28429), .S(n29462), .Y(n28436) );
  MUX2X1 U18768 ( .B(n28435), .A(n28420), .S(n28609), .Y(n28469) );
  MUX2X1 U18769 ( .B(grid[183]), .A(grid[189]), .S(n26153), .Y(n28440) );
  MUX2X1 U18770 ( .B(grid[171]), .A(grid[177]), .S(n26086), .Y(n28439) );
  MUX2X1 U18771 ( .B(grid[159]), .A(grid[165]), .S(n26123), .Y(n28443) );
  MUX2X1 U18772 ( .B(grid[147]), .A(grid[153]), .S(n26109), .Y(n28442) );
  MUX2X1 U18773 ( .B(n28441), .A(n28438), .S(n26304), .Y(n28452) );
  MUX2X1 U18774 ( .B(grid[135]), .A(grid[141]), .S(n26153), .Y(n28446) );
  MUX2X1 U18775 ( .B(grid[123]), .A(grid[129]), .S(n26103), .Y(n28445) );
  MUX2X1 U18776 ( .B(grid[111]), .A(grid[117]), .S(n26087), .Y(n28449) );
  MUX2X1 U18777 ( .B(grid[99]), .A(grid[105]), .S(n26088), .Y(n28448) );
  MUX2X1 U18778 ( .B(n28447), .A(n28444), .S(n29462), .Y(n28451) );
  MUX2X1 U18779 ( .B(grid[87]), .A(grid[93]), .S(n26144), .Y(n28455) );
  MUX2X1 U18780 ( .B(grid[75]), .A(grid[81]), .S(n26120), .Y(n28454) );
  MUX2X1 U18781 ( .B(grid[63]), .A(grid[69]), .S(n26143), .Y(n28458) );
  MUX2X1 U18782 ( .B(grid[51]), .A(grid[57]), .S(n26079), .Y(n28457) );
  MUX2X1 U18783 ( .B(n28456), .A(n28453), .S(n29462), .Y(n28467) );
  MUX2X1 U18784 ( .B(grid[39]), .A(grid[45]), .S(n26113), .Y(n28461) );
  MUX2X1 U18785 ( .B(grid[27]), .A(grid[33]), .S(n26093), .Y(n28460) );
  MUX2X1 U18786 ( .B(grid[15]), .A(grid[21]), .S(n26084), .Y(n28464) );
  MUX2X1 U18787 ( .B(grid[3]), .A(grid[9]), .S(n26115), .Y(n28463) );
  MUX2X1 U18788 ( .B(n28462), .A(n28459), .S(n29462), .Y(n28466) );
  MUX2X1 U18789 ( .B(n28465), .A(n28450), .S(n28609), .Y(n28468) );
  MUX2X1 U18790 ( .B(grid[376]), .A(grid[382]), .S(n26119), .Y(n28472) );
  MUX2X1 U18791 ( .B(grid[364]), .A(grid[370]), .S(n26112), .Y(n28471) );
  MUX2X1 U18792 ( .B(grid[352]), .A(grid[358]), .S(n26090), .Y(n28475) );
  MUX2X1 U18793 ( .B(grid[340]), .A(grid[346]), .S(n26107), .Y(n28474) );
  MUX2X1 U18794 ( .B(n28473), .A(n28470), .S(n26304), .Y(n28484) );
  MUX2X1 U18795 ( .B(grid[328]), .A(grid[334]), .S(n26146), .Y(n28478) );
  MUX2X1 U18796 ( .B(grid[304]), .A(grid[310]), .S(n26141), .Y(n28481) );
  MUX2X1 U18797 ( .B(grid[292]), .A(grid[298]), .S(n26143), .Y(n28480) );
  MUX2X1 U18798 ( .B(n28479), .A(n28476), .S(n29462), .Y(n28483) );
  MUX2X1 U18799 ( .B(grid[280]), .A(grid[286]), .S(n26140), .Y(n28487) );
  MUX2X1 U18800 ( .B(grid[268]), .A(grid[274]), .S(n26095), .Y(n28486) );
  MUX2X1 U18801 ( .B(grid[256]), .A(grid[262]), .S(n26121), .Y(n28490) );
  MUX2X1 U18802 ( .B(grid[244]), .A(grid[250]), .S(n26122), .Y(n28489) );
  MUX2X1 U18803 ( .B(n28488), .A(n28485), .S(n21129), .Y(n28499) );
  MUX2X1 U18804 ( .B(grid[232]), .A(grid[238]), .S(n26120), .Y(n28493) );
  MUX2X1 U18805 ( .B(grid[220]), .A(grid[226]), .S(n26144), .Y(n28492) );
  MUX2X1 U18806 ( .B(grid[208]), .A(grid[214]), .S(n26102), .Y(n28496) );
  MUX2X1 U18807 ( .B(grid[196]), .A(grid[202]), .S(n26128), .Y(n28495) );
  MUX2X1 U18808 ( .B(n28494), .A(n28491), .S(n21129), .Y(n28498) );
  MUX2X1 U18809 ( .B(n28497), .A(n28482), .S(n28609), .Y(n28531) );
  MUX2X1 U18810 ( .B(grid[184]), .A(grid[190]), .S(n26096), .Y(n28502) );
  MUX2X1 U18811 ( .B(grid[160]), .A(grid[166]), .S(n26089), .Y(n28505) );
  MUX2X1 U18812 ( .B(grid[148]), .A(grid[154]), .S(n26149), .Y(n28504) );
  MUX2X1 U18813 ( .B(grid[136]), .A(grid[142]), .S(n26134), .Y(n28508) );
  MUX2X1 U18814 ( .B(grid[112]), .A(grid[118]), .S(n26089), .Y(n28511) );
  MUX2X1 U18815 ( .B(n28509), .A(n28506), .S(n21129), .Y(n28513) );
  MUX2X1 U18816 ( .B(grid[88]), .A(grid[94]), .S(n25592), .Y(n28517) );
  MUX2X1 U18817 ( .B(grid[76]), .A(grid[82]), .S(n26150), .Y(n28516) );
  MUX2X1 U18818 ( .B(grid[64]), .A(grid[70]), .S(n26135), .Y(n28520) );
  MUX2X1 U18819 ( .B(grid[40]), .A(grid[46]), .S(n26151), .Y(n28523) );
  MUX2X1 U18820 ( .B(grid[28]), .A(grid[34]), .S(n23208), .Y(n28522) );
  MUX2X1 U18821 ( .B(grid[16]), .A(grid[22]), .S(n26139), .Y(n28526) );
  MUX2X1 U18822 ( .B(n28527), .A(n28512), .S(n28609), .Y(n28530) );
  MUX2X1 U18823 ( .B(grid[377]), .A(grid[383]), .S(n26085), .Y(n28534) );
  MUX2X1 U18824 ( .B(grid[365]), .A(grid[371]), .S(n26124), .Y(n28533) );
  MUX2X1 U18825 ( .B(grid[353]), .A(grid[359]), .S(n26090), .Y(n28537) );
  MUX2X1 U18826 ( .B(grid[341]), .A(grid[347]), .S(n26111), .Y(n28536) );
  MUX2X1 U18827 ( .B(n28535), .A(n28532), .S(n26304), .Y(n28546) );
  MUX2X1 U18828 ( .B(grid[329]), .A(grid[335]), .S(n26125), .Y(n28540) );
  MUX2X1 U18829 ( .B(grid[317]), .A(grid[323]), .S(n26097), .Y(n28539) );
  MUX2X1 U18830 ( .B(grid[305]), .A(grid[311]), .S(n26103), .Y(n28543) );
  MUX2X1 U18831 ( .B(grid[293]), .A(grid[299]), .S(n26082), .Y(n28542) );
  MUX2X1 U18832 ( .B(n28541), .A(n28538), .S(n29462), .Y(n28545) );
  MUX2X1 U18833 ( .B(grid[281]), .A(grid[287]), .S(n26142), .Y(n28549) );
  MUX2X1 U18834 ( .B(grid[269]), .A(grid[275]), .S(n26095), .Y(n28548) );
  MUX2X1 U18835 ( .B(grid[257]), .A(grid[263]), .S(n26094), .Y(n28552) );
  MUX2X1 U18836 ( .B(grid[245]), .A(grid[251]), .S(n26112), .Y(n28551) );
  MUX2X1 U18837 ( .B(n28550), .A(n28547), .S(n21129), .Y(n28561) );
  MUX2X1 U18838 ( .B(grid[233]), .A(grid[239]), .S(n26106), .Y(n28555) );
  MUX2X1 U18839 ( .B(grid[221]), .A(grid[227]), .S(n26088), .Y(n28554) );
  MUX2X1 U18840 ( .B(grid[209]), .A(grid[215]), .S(n26117), .Y(n28558) );
  MUX2X1 U18841 ( .B(grid[197]), .A(grid[203]), .S(n26141), .Y(n28557) );
  MUX2X1 U18842 ( .B(n28559), .A(n28544), .S(n28609), .Y(n28593) );
  MUX2X1 U18843 ( .B(grid[185]), .A(grid[191]), .S(n26094), .Y(n28564) );
  MUX2X1 U18844 ( .B(grid[161]), .A(grid[167]), .S(n26097), .Y(n28567) );
  MUX2X1 U18845 ( .B(grid[149]), .A(grid[155]), .S(n26148), .Y(n28566) );
  MUX2X1 U18846 ( .B(n28565), .A(n28562), .S(n29462), .Y(n28576) );
  MUX2X1 U18847 ( .B(grid[125]), .A(grid[131]), .S(n26093), .Y(n28569) );
  MUX2X1 U18848 ( .B(grid[113]), .A(grid[119]), .S(n26137), .Y(n28573) );
  MUX2X1 U18849 ( .B(grid[101]), .A(grid[107]), .S(n26101), .Y(n28572) );
  MUX2X1 U18850 ( .B(n28571), .A(n28568), .S(n21129), .Y(n28575) );
  MUX2X1 U18851 ( .B(grid[89]), .A(grid[95]), .S(n26108), .Y(n28579) );
  MUX2X1 U18852 ( .B(grid[77]), .A(grid[83]), .S(n25592), .Y(n28578) );
  MUX2X1 U18853 ( .B(grid[65]), .A(grid[71]), .S(n26125), .Y(n28582) );
  MUX2X1 U18854 ( .B(grid[53]), .A(grid[59]), .S(n26153), .Y(n28581) );
  MUX2X1 U18855 ( .B(grid[41]), .A(grid[47]), .S(n26145), .Y(n28585) );
  MUX2X1 U18856 ( .B(grid[29]), .A(grid[35]), .S(n26130), .Y(n28584) );
  MUX2X1 U18857 ( .B(grid[17]), .A(grid[23]), .S(n26146), .Y(n28588) );
  MUX2X1 U18858 ( .B(n28586), .A(n28583), .S(n21129), .Y(n28590) );
  MUX2X1 U18859 ( .B(n28589), .A(n28574), .S(n28609), .Y(n28592) );
  MUX2X1 U18860 ( .B(n28611), .A(n28612), .S(n26398), .Y(n28610) );
  MUX2X1 U18861 ( .B(n28614), .A(n28615), .S(n26428), .Y(n28613) );
  MUX2X1 U18862 ( .B(n28617), .A(n28618), .S(n26349), .Y(n28616) );
  MUX2X1 U18863 ( .B(n28620), .A(n28621), .S(n26352), .Y(n28619) );
  MUX2X1 U18864 ( .B(n28623), .A(n28624), .S(n27214), .Y(n28622) );
  MUX2X1 U18865 ( .B(n28626), .A(n28627), .S(n26427), .Y(n28625) );
  MUX2X1 U18866 ( .B(n28629), .A(n28630), .S(n26430), .Y(n28628) );
  MUX2X1 U18867 ( .B(n28632), .A(n28633), .S(n26351), .Y(n28631) );
  MUX2X1 U18868 ( .B(n28635), .A(n28636), .S(n26396), .Y(n28634) );
  MUX2X1 U18869 ( .B(n28638), .A(n28639), .S(n27214), .Y(n28637) );
  MUX2X1 U18870 ( .B(n28641), .A(n28642), .S(n26348), .Y(n28640) );
  MUX2X1 U18871 ( .B(n28644), .A(n28645), .S(n26350), .Y(n28643) );
  MUX2X1 U18872 ( .B(n28647), .A(n28648), .S(n26412), .Y(n28646) );
  MUX2X1 U18873 ( .B(n28650), .A(n28651), .S(n26418), .Y(n28649) );
  MUX2X1 U18874 ( .B(n28653), .A(n28654), .S(n27214), .Y(n28652) );
  MUX2X1 U18875 ( .B(n28656), .A(n28657), .S(n26378), .Y(n28655) );
  MUX2X1 U18876 ( .B(n28659), .A(n28660), .S(n26397), .Y(n28658) );
  MUX2X1 U18877 ( .B(n28662), .A(n28663), .S(n26419), .Y(n28661) );
  MUX2X1 U18878 ( .B(n28665), .A(n28666), .S(n26355), .Y(n28664) );
  MUX2X1 U18879 ( .B(n28668), .A(n28669), .S(n27214), .Y(n28667) );
  MUX2X1 U18880 ( .B(n28670), .A(n28671), .S(n26481), .Y(n13804) );
  MUX2X1 U18881 ( .B(n28673), .A(n28674), .S(n26434), .Y(n28672) );
  MUX2X1 U18882 ( .B(n28676), .A(n28677), .S(n26436), .Y(n28675) );
  MUX2X1 U18883 ( .B(n28679), .A(n28680), .S(n26399), .Y(n28678) );
  MUX2X1 U18884 ( .B(n28682), .A(n28683), .S(n26429), .Y(n28681) );
  MUX2X1 U18885 ( .B(n28685), .A(n28686), .S(n27214), .Y(n28684) );
  MUX2X1 U18886 ( .B(n28688), .A(n28689), .S(n26435), .Y(n28687) );
  MUX2X1 U18887 ( .B(n28691), .A(n28692), .S(n26437), .Y(n28690) );
  MUX2X1 U18888 ( .B(n28694), .A(n28695), .S(n26370), .Y(n28693) );
  MUX2X1 U18889 ( .B(n28697), .A(n28698), .S(n26431), .Y(n28696) );
  MUX2X1 U18890 ( .B(n28700), .A(n28701), .S(n27214), .Y(n28699) );
  MUX2X1 U18891 ( .B(n28703), .A(n28704), .S(n26438), .Y(n28702) );
  MUX2X1 U18892 ( .B(n28706), .A(n28707), .S(n26440), .Y(n28705) );
  MUX2X1 U18893 ( .B(n28709), .A(n28710), .S(n26432), .Y(n28708) );
  MUX2X1 U18894 ( .B(n28712), .A(n28713), .S(n26433), .Y(n28711) );
  MUX2X1 U18895 ( .B(n28715), .A(n28716), .S(n27214), .Y(n28714) );
  MUX2X1 U18896 ( .B(n28718), .A(n28719), .S(n26439), .Y(n28717) );
  MUX2X1 U18897 ( .B(n28721), .A(n28722), .S(n26442), .Y(n28720) );
  MUX2X1 U18898 ( .B(n28724), .A(n28725), .S(n26367), .Y(n28723) );
  MUX2X1 U18899 ( .B(n28727), .A(n28728), .S(n26443), .Y(n28726) );
  MUX2X1 U18900 ( .B(n28730), .A(n28731), .S(n27214), .Y(n28729) );
  MUX2X1 U18901 ( .B(n28732), .A(n28733), .S(n26481), .Y(n13803) );
  MUX2X1 U18902 ( .B(n28735), .A(n28736), .S(n26379), .Y(n28734) );
  MUX2X1 U18903 ( .B(n28738), .A(n28739), .S(n26383), .Y(n28737) );
  MUX2X1 U18904 ( .B(n28741), .A(n28742), .S(n26421), .Y(n28740) );
  MUX2X1 U18905 ( .B(n28744), .A(n28745), .S(n26361), .Y(n28743) );
  MUX2X1 U18906 ( .B(n28747), .A(n28748), .S(n27214), .Y(n28746) );
  MUX2X1 U18907 ( .B(n28750), .A(n28751), .S(n26417), .Y(n28749) );
  MUX2X1 U18908 ( .B(n28753), .A(n28754), .S(n26356), .Y(n28752) );
  MUX2X1 U18909 ( .B(n28756), .A(n28757), .S(n26422), .Y(n28755) );
  MUX2X1 U18910 ( .B(n28759), .A(n28760), .S(n26362), .Y(n28758) );
  MUX2X1 U18911 ( .B(n28762), .A(n28763), .S(n27214), .Y(n28761) );
  MUX2X1 U18912 ( .B(n28765), .A(n28766), .S(n26420), .Y(n28764) );
  MUX2X1 U18913 ( .B(n28768), .A(n28769), .S(n26359), .Y(n28767) );
  MUX2X1 U18914 ( .B(n28771), .A(n28772), .S(n26406), .Y(n28770) );
  MUX2X1 U18915 ( .B(n28774), .A(n28775), .S(n26414), .Y(n28773) );
  MUX2X1 U18916 ( .B(n28777), .A(n28778), .S(n27214), .Y(n28776) );
  MUX2X1 U18917 ( .B(n28780), .A(n28781), .S(n26358), .Y(n28779) );
  MUX2X1 U18918 ( .B(n28783), .A(n28784), .S(n26343), .Y(n28782) );
  MUX2X1 U18919 ( .B(n28786), .A(n28787), .S(n26413), .Y(n28785) );
  MUX2X1 U18920 ( .B(n28789), .A(n28790), .S(n26383), .Y(n28788) );
  MUX2X1 U18921 ( .B(n28792), .A(n28793), .S(n27214), .Y(n28791) );
  MUX2X1 U18922 ( .B(n28794), .A(n28795), .S(n26482), .Y(n13802) );
  MUX2X1 U18923 ( .B(n28797), .A(n28798), .S(n26371), .Y(n28796) );
  MUX2X1 U18924 ( .B(n28800), .A(n28801), .S(n26386), .Y(n28799) );
  MUX2X1 U18925 ( .B(n28803), .A(n28804), .S(n26374), .Y(n28802) );
  MUX2X1 U18926 ( .B(n28806), .A(n28807), .S(n26394), .Y(n28805) );
  MUX2X1 U18927 ( .B(n28809), .A(n28810), .S(n27214), .Y(n28808) );
  MUX2X1 U18928 ( .B(n28812), .A(n28813), .S(n26385), .Y(n28811) );
  MUX2X1 U18929 ( .B(n28815), .A(n28816), .S(n26441), .Y(n28814) );
  MUX2X1 U18930 ( .B(n28818), .A(n28819), .S(n26391), .Y(n28817) );
  MUX2X1 U18931 ( .B(n28821), .A(n28822), .S(n26372), .Y(n28820) );
  MUX2X1 U18932 ( .B(n28824), .A(n28825), .S(n27214), .Y(n28823) );
  MUX2X1 U18933 ( .B(n28827), .A(n28828), .S(n26374), .Y(n28826) );
  MUX2X1 U18934 ( .B(n28830), .A(n28831), .S(n26393), .Y(n28829) );
  MUX2X1 U18935 ( .B(n28833), .A(n28834), .S(n26390), .Y(n28832) );
  MUX2X1 U18936 ( .B(n28836), .A(n28837), .S(n26368), .Y(n28835) );
  MUX2X1 U18937 ( .B(n28839), .A(n28840), .S(n27214), .Y(n28838) );
  MUX2X1 U18938 ( .B(n28842), .A(n28843), .S(n26392), .Y(n28841) );
  MUX2X1 U18939 ( .B(n28845), .A(n28846), .S(n26443), .Y(n28844) );
  MUX2X1 U18940 ( .B(n28848), .A(n28849), .S(n26369), .Y(n28847) );
  MUX2X1 U18941 ( .B(n28851), .A(n28852), .S(n26384), .Y(n28850) );
  MUX2X1 U18942 ( .B(n28854), .A(n28855), .S(n27214), .Y(n28853) );
  MUX2X1 U18943 ( .B(n28856), .A(n28857), .S(n26482), .Y(n13801) );
  MUX2X1 U18944 ( .B(n28859), .A(n28860), .S(n26415), .Y(n28858) );
  MUX2X1 U18945 ( .B(n28862), .A(n28863), .S(n26373), .Y(n28861) );
  MUX2X1 U18946 ( .B(n28865), .A(n28866), .S(n26373), .Y(n28864) );
  MUX2X1 U18947 ( .B(n28868), .A(n28869), .S(n26408), .Y(n28867) );
  MUX2X1 U18948 ( .B(n28871), .A(n28872), .S(n27214), .Y(n28870) );
  MUX2X1 U18949 ( .B(n28874), .A(n28875), .S(n26372), .Y(n28873) );
  MUX2X1 U18950 ( .B(n28877), .A(n28878), .S(n26387), .Y(n28876) );
  MUX2X1 U18951 ( .B(n28880), .A(n28881), .S(n26407), .Y(n28879) );
  MUX2X1 U18952 ( .B(n28883), .A(n28884), .S(n26395), .Y(n28882) );
  MUX2X1 U18953 ( .B(n28886), .A(n28887), .S(n27214), .Y(n28885) );
  MUX2X1 U18954 ( .B(n28889), .A(n28890), .S(n26416), .Y(n28888) );
  MUX2X1 U18955 ( .B(n28892), .A(n28893), .S(n26409), .Y(n28891) );
  MUX2X1 U18956 ( .B(n28895), .A(n28896), .S(n26375), .Y(n28894) );
  MUX2X1 U18957 ( .B(n28898), .A(n28899), .S(n26410), .Y(n28897) );
  MUX2X1 U18958 ( .B(n28901), .A(n28902), .S(n27214), .Y(n28900) );
  MUX2X1 U18959 ( .B(n28904), .A(n28905), .S(n26375), .Y(n28903) );
  MUX2X1 U18960 ( .B(n28907), .A(n28908), .S(n26367), .Y(n28906) );
  MUX2X1 U18961 ( .B(n28910), .A(n28911), .S(n26371), .Y(n28909) );
  MUX2X1 U18962 ( .B(n28913), .A(n28914), .S(n26370), .Y(n28912) );
  MUX2X1 U18963 ( .B(n28916), .A(n28917), .S(n27214), .Y(n28915) );
  MUX2X1 U18964 ( .B(n28918), .A(n28919), .S(n26483), .Y(n13800) );
  MUX2X1 U18965 ( .B(n28921), .A(n28922), .S(n26380), .Y(n28920) );
  MUX2X1 U18966 ( .B(n28924), .A(n28925), .S(n26382), .Y(n28923) );
  MUX2X1 U18967 ( .B(n28927), .A(n28928), .S(n26380), .Y(n28926) );
  MUX2X1 U18968 ( .B(n28930), .A(n28931), .S(n26364), .Y(n28929) );
  MUX2X1 U18969 ( .B(n28933), .A(n28934), .S(n27214), .Y(n28932) );
  MUX2X1 U18970 ( .B(n28936), .A(n28937), .S(n26381), .Y(n28935) );
  MUX2X1 U18971 ( .B(n28939), .A(n28940), .S(n26360), .Y(n28938) );
  MUX2X1 U18972 ( .B(n28942), .A(n28943), .S(n26363), .Y(n28941) );
  MUX2X1 U18973 ( .B(n28945), .A(n28946), .S(n26347), .Y(n28944) );
  MUX2X1 U18974 ( .B(n28948), .A(n28949), .S(n27214), .Y(n28947) );
  MUX2X1 U18975 ( .B(n28951), .A(n28952), .S(n26357), .Y(n28950) );
  MUX2X1 U18976 ( .B(n28954), .A(n28955), .S(n26345), .Y(n28953) );
  MUX2X1 U18977 ( .B(n28957), .A(n28958), .S(n26405), .Y(n28956) );
  MUX2X1 U18978 ( .B(n28960), .A(n28961), .S(n26411), .Y(n28959) );
  MUX2X1 U18979 ( .B(n28963), .A(n28964), .S(n27214), .Y(n28962) );
  MUX2X1 U18980 ( .B(n28966), .A(n28967), .S(n26344), .Y(n28965) );
  MUX2X1 U18981 ( .B(n28969), .A(n28970), .S(n26346), .Y(n28968) );
  MUX2X1 U18982 ( .B(n28972), .A(n28973), .S(n26382), .Y(n28971) );
  MUX2X1 U18983 ( .B(n28975), .A(n28976), .S(n26379), .Y(n28974) );
  MUX2X1 U18984 ( .B(n28978), .A(n28979), .S(n27214), .Y(n28977) );
  MUX2X1 U18985 ( .B(n28980), .A(n28981), .S(n26483), .Y(n13799) );
  MUX2X1 U18986 ( .B(grid[372]), .A(grid[378]), .S(n26177), .Y(n28612) );
  MUX2X1 U18987 ( .B(grid[360]), .A(grid[366]), .S(n26188), .Y(n28611) );
  MUX2X1 U18988 ( .B(grid[348]), .A(grid[354]), .S(n26226), .Y(n28615) );
  MUX2X1 U18989 ( .B(grid[336]), .A(grid[342]), .S(n26214), .Y(n28614) );
  MUX2X1 U18990 ( .B(n28613), .A(n28610), .S(n26543), .Y(n28624) );
  MUX2X1 U18991 ( .B(grid[324]), .A(grid[330]), .S(n26187), .Y(n28618) );
  MUX2X1 U18992 ( .B(grid[312]), .A(grid[318]), .S(n26186), .Y(n28617) );
  MUX2X1 U18993 ( .B(grid[300]), .A(grid[306]), .S(n26213), .Y(n28621) );
  MUX2X1 U18994 ( .B(grid[288]), .A(grid[294]), .S(n26224), .Y(n28620) );
  MUX2X1 U18995 ( .B(n28619), .A(n28616), .S(n26568), .Y(n28623) );
  MUX2X1 U18996 ( .B(grid[276]), .A(grid[282]), .S(n26227), .Y(n28627) );
  MUX2X1 U18997 ( .B(grid[264]), .A(grid[270]), .S(n26262), .Y(n28626) );
  MUX2X1 U18998 ( .B(grid[252]), .A(grid[258]), .S(n26199), .Y(n28630) );
  MUX2X1 U18999 ( .B(grid[240]), .A(grid[246]), .S(n26173), .Y(n28629) );
  MUX2X1 U19000 ( .B(n28628), .A(n28625), .S(n26527), .Y(n28639) );
  MUX2X1 U19001 ( .B(grid[228]), .A(grid[234]), .S(n26212), .Y(n28633) );
  MUX2X1 U19002 ( .B(grid[216]), .A(grid[222]), .S(n26176), .Y(n28632) );
  MUX2X1 U19003 ( .B(grid[192]), .A(grid[198]), .S(n26182), .Y(n28635) );
  MUX2X1 U19004 ( .B(n28634), .A(n28631), .S(n26571), .Y(n28638) );
  MUX2X1 U19005 ( .B(n28637), .A(n28622), .S(n28993), .Y(n28671) );
  MUX2X1 U19006 ( .B(grid[180]), .A(grid[186]), .S(n26186), .Y(n28642) );
  MUX2X1 U19007 ( .B(grid[168]), .A(grid[174]), .S(n26185), .Y(n28641) );
  MUX2X1 U19008 ( .B(grid[156]), .A(grid[162]), .S(n26211), .Y(n28645) );
  MUX2X1 U19009 ( .B(grid[144]), .A(grid[150]), .S(n26175), .Y(n28644) );
  MUX2X1 U19010 ( .B(n28643), .A(n28640), .S(n26567), .Y(n28654) );
  MUX2X1 U19011 ( .B(grid[132]), .A(grid[138]), .S(n26184), .Y(n28648) );
  MUX2X1 U19012 ( .B(grid[120]), .A(grid[126]), .S(n26198), .Y(n28647) );
  MUX2X1 U19013 ( .B(grid[108]), .A(grid[114]), .S(n26174), .Y(n28651) );
  MUX2X1 U19014 ( .B(grid[96]), .A(grid[102]), .S(n26214), .Y(n28650) );
  MUX2X1 U19015 ( .B(n28649), .A(n28646), .S(n26562), .Y(n28653) );
  MUX2X1 U19016 ( .B(grid[84]), .A(grid[90]), .S(n26261), .Y(n28657) );
  MUX2X1 U19017 ( .B(grid[72]), .A(grid[78]), .S(n26178), .Y(n28656) );
  MUX2X1 U19018 ( .B(grid[60]), .A(grid[66]), .S(n26172), .Y(n28660) );
  MUX2X1 U19019 ( .B(grid[48]), .A(grid[54]), .S(n26183), .Y(n28659) );
  MUX2X1 U19020 ( .B(n28658), .A(n28655), .S(n26569), .Y(n28669) );
  MUX2X1 U19021 ( .B(grid[36]), .A(grid[42]), .S(n26177), .Y(n28663) );
  MUX2X1 U19022 ( .B(grid[24]), .A(grid[30]), .S(n26215), .Y(n28662) );
  MUX2X1 U19023 ( .B(grid[12]), .A(grid[18]), .S(n26184), .Y(n28666) );
  MUX2X1 U19024 ( .B(grid[0]), .A(grid[6]), .S(n26244), .Y(n28665) );
  MUX2X1 U19025 ( .B(n28664), .A(n28661), .S(n26563), .Y(n28668) );
  MUX2X1 U19026 ( .B(n28667), .A(n28652), .S(n28993), .Y(n28670) );
  MUX2X1 U19027 ( .B(grid[373]), .A(grid[379]), .S(n26196), .Y(n28674) );
  MUX2X1 U19028 ( .B(grid[361]), .A(grid[367]), .S(n26225), .Y(n28673) );
  MUX2X1 U19029 ( .B(grid[349]), .A(grid[355]), .S(n26197), .Y(n28677) );
  MUX2X1 U19030 ( .B(grid[337]), .A(grid[343]), .S(n26197), .Y(n28676) );
  MUX2X1 U19031 ( .B(n28675), .A(n28672), .S(n26534), .Y(n28686) );
  MUX2X1 U19032 ( .B(grid[325]), .A(grid[331]), .S(n26178), .Y(n28680) );
  MUX2X1 U19033 ( .B(grid[313]), .A(grid[319]), .S(n26202), .Y(n28679) );
  MUX2X1 U19034 ( .B(grid[301]), .A(grid[307]), .S(n26228), .Y(n28683) );
  MUX2X1 U19035 ( .B(grid[289]), .A(grid[295]), .S(n26264), .Y(n28682) );
  MUX2X1 U19036 ( .B(n28681), .A(n28678), .S(n26525), .Y(n28685) );
  MUX2X1 U19037 ( .B(grid[277]), .A(grid[283]), .S(n26198), .Y(n28689) );
  MUX2X1 U19038 ( .B(grid[265]), .A(grid[271]), .S(n26198), .Y(n28688) );
  MUX2X1 U19039 ( .B(grid[253]), .A(grid[259]), .S(n26199), .Y(n28692) );
  MUX2X1 U19040 ( .B(grid[241]), .A(grid[247]), .S(n26230), .Y(n28691) );
  MUX2X1 U19041 ( .B(grid[229]), .A(grid[235]), .S(n26229), .Y(n28695) );
  MUX2X1 U19042 ( .B(grid[217]), .A(grid[223]), .S(n26265), .Y(n28694) );
  MUX2X1 U19043 ( .B(grid[205]), .A(grid[211]), .S(n26229), .Y(n28698) );
  MUX2X1 U19044 ( .B(grid[193]), .A(grid[199]), .S(n26175), .Y(n28697) );
  MUX2X1 U19045 ( .B(n28696), .A(n28693), .S(n26530), .Y(n28700) );
  MUX2X1 U19046 ( .B(n28699), .A(n28684), .S(n28993), .Y(n28733) );
  MUX2X1 U19047 ( .B(grid[181]), .A(grid[187]), .S(n26224), .Y(n28704) );
  MUX2X1 U19048 ( .B(grid[169]), .A(grid[175]), .S(n26210), .Y(n28703) );
  MUX2X1 U19049 ( .B(grid[157]), .A(grid[163]), .S(n26230), .Y(n28707) );
  MUX2X1 U19050 ( .B(grid[145]), .A(grid[151]), .S(n26266), .Y(n28706) );
  MUX2X1 U19051 ( .B(n28705), .A(n28702), .S(n26576), .Y(n28716) );
  MUX2X1 U19052 ( .B(grid[133]), .A(grid[139]), .S(n26201), .Y(n28710) );
  MUX2X1 U19053 ( .B(grid[121]), .A(grid[127]), .S(n26173), .Y(n28709) );
  MUX2X1 U19054 ( .B(grid[109]), .A(grid[115]), .S(n26263), .Y(n28713) );
  MUX2X1 U19055 ( .B(grid[97]), .A(grid[103]), .S(n26226), .Y(n28712) );
  MUX2X1 U19056 ( .B(n28711), .A(n28708), .S(n26553), .Y(n28715) );
  MUX2X1 U19057 ( .B(grid[85]), .A(grid[91]), .S(n26196), .Y(n28719) );
  MUX2X1 U19058 ( .B(grid[73]), .A(grid[79]), .S(n26267), .Y(n28718) );
  MUX2X1 U19059 ( .B(grid[61]), .A(grid[67]), .S(n26200), .Y(n28722) );
  MUX2X1 U19060 ( .B(grid[49]), .A(grid[55]), .S(n26176), .Y(n28721) );
  MUX2X1 U19061 ( .B(n28720), .A(n28717), .S(n26570), .Y(n28731) );
  MUX2X1 U19062 ( .B(n25480), .A(grid[43]), .S(n26262), .Y(n28725) );
  MUX2X1 U19063 ( .B(grid[25]), .A(grid[31]), .S(n26225), .Y(n28724) );
  MUX2X1 U19064 ( .B(grid[13]), .A(grid[19]), .S(n26174), .Y(n28728) );
  MUX2X1 U19065 ( .B(grid[1]), .A(grid[7]), .S(n26185), .Y(n28727) );
  MUX2X1 U19066 ( .B(n28726), .A(n28723), .S(n26558), .Y(n28730) );
  MUX2X1 U19067 ( .B(n28729), .A(n28714), .S(n28993), .Y(n28732) );
  MUX2X1 U19068 ( .B(grid[374]), .A(grid[380]), .S(n26252), .Y(n28736) );
  MUX2X1 U19069 ( .B(grid[362]), .A(grid[368]), .S(n26182), .Y(n28735) );
  MUX2X1 U19070 ( .B(grid[350]), .A(grid[356]), .S(n26187), .Y(n28739) );
  MUX2X1 U19071 ( .B(grid[338]), .A(grid[344]), .S(n26267), .Y(n28738) );
  MUX2X1 U19072 ( .B(n28737), .A(n28734), .S(n26574), .Y(n28748) );
  MUX2X1 U19073 ( .B(grid[326]), .A(grid[332]), .S(n26258), .Y(n28742) );
  MUX2X1 U19074 ( .B(grid[314]), .A(grid[320]), .S(n26256), .Y(n28741) );
  MUX2X1 U19075 ( .B(grid[302]), .A(grid[308]), .S(n26266), .Y(n28745) );
  MUX2X1 U19076 ( .B(n25610), .A(grid[296]), .S(n26265), .Y(n28744) );
  MUX2X1 U19077 ( .B(n28743), .A(n28740), .S(n26545), .Y(n28747) );
  MUX2X1 U19078 ( .B(n25465), .A(grid[284]), .S(n26188), .Y(n28751) );
  MUX2X1 U19079 ( .B(grid[266]), .A(grid[272]), .S(n26268), .Y(n28750) );
  MUX2X1 U19080 ( .B(grid[254]), .A(grid[260]), .S(n26185), .Y(n28754) );
  MUX2X1 U19081 ( .B(grid[242]), .A(grid[248]), .S(n26238), .Y(n28753) );
  MUX2X1 U19082 ( .B(n28752), .A(n28749), .S(n26575), .Y(n28763) );
  MUX2X1 U19083 ( .B(grid[230]), .A(grid[236]), .S(n26199), .Y(n28757) );
  MUX2X1 U19084 ( .B(grid[218]), .A(grid[224]), .S(n26266), .Y(n28756) );
  MUX2X1 U19085 ( .B(grid[206]), .A(grid[212]), .S(n26216), .Y(n28760) );
  MUX2X1 U19086 ( .B(n25505), .A(grid[200]), .S(n26252), .Y(n28759) );
  MUX2X1 U19087 ( .B(n28758), .A(n28755), .S(n26528), .Y(n28762) );
  MUX2X1 U19088 ( .B(n28761), .A(n28746), .S(n28993), .Y(n28795) );
  MUX2X1 U19089 ( .B(grid[182]), .A(grid[188]), .S(n26183), .Y(n28766) );
  MUX2X1 U19090 ( .B(grid[170]), .A(grid[176]), .S(n26258), .Y(n28765) );
  MUX2X1 U19091 ( .B(grid[158]), .A(grid[164]), .S(n26200), .Y(n28769) );
  MUX2X1 U19092 ( .B(grid[146]), .A(grid[152]), .S(n26173), .Y(n28768) );
  MUX2X1 U19093 ( .B(n28767), .A(n28764), .S(n26546), .Y(n28778) );
  MUX2X1 U19094 ( .B(grid[134]), .A(grid[140]), .S(n26257), .Y(n28772) );
  MUX2X1 U19095 ( .B(grid[122]), .A(grid[128]), .S(n26215), .Y(n28771) );
  MUX2X1 U19096 ( .B(grid[110]), .A(grid[116]), .S(n26267), .Y(n28775) );
  MUX2X1 U19097 ( .B(grid[98]), .A(grid[104]), .S(n26178), .Y(n28774) );
  MUX2X1 U19098 ( .B(n28773), .A(n28770), .S(n26544), .Y(n28777) );
  MUX2X1 U19099 ( .B(grid[86]), .A(grid[92]), .S(n26172), .Y(n28781) );
  MUX2X1 U19100 ( .B(grid[74]), .A(grid[80]), .S(n26172), .Y(n28780) );
  MUX2X1 U19101 ( .B(grid[62]), .A(grid[68]), .S(n26239), .Y(n28784) );
  MUX2X1 U19102 ( .B(grid[50]), .A(grid[56]), .S(n26244), .Y(n28783) );
  MUX2X1 U19103 ( .B(n28782), .A(n28779), .S(n26529), .Y(n28793) );
  MUX2X1 U19104 ( .B(grid[38]), .A(grid[44]), .S(n26268), .Y(n28787) );
  MUX2X1 U19105 ( .B(grid[26]), .A(grid[32]), .S(n26224), .Y(n28786) );
  MUX2X1 U19106 ( .B(grid[14]), .A(grid[20]), .S(n26243), .Y(n28790) );
  MUX2X1 U19107 ( .B(grid[2]), .A(grid[8]), .S(n26201), .Y(n28789) );
  MUX2X1 U19108 ( .B(n28788), .A(n28785), .S(n26546), .Y(n28792) );
  MUX2X1 U19109 ( .B(n28791), .A(n28776), .S(n28993), .Y(n28794) );
  MUX2X1 U19110 ( .B(grid[375]), .A(grid[381]), .S(n26255), .Y(n28798) );
  MUX2X1 U19111 ( .B(grid[363]), .A(grid[369]), .S(n26254), .Y(n28797) );
  MUX2X1 U19112 ( .B(grid[351]), .A(grid[357]), .S(n26175), .Y(n28801) );
  MUX2X1 U19113 ( .B(grid[339]), .A(grid[345]), .S(n26262), .Y(n28800) );
  MUX2X1 U19114 ( .B(n28799), .A(n28796), .S(n26564), .Y(n28810) );
  MUX2X1 U19115 ( .B(grid[327]), .A(grid[333]), .S(n26243), .Y(n28804) );
  MUX2X1 U19116 ( .B(grid[315]), .A(grid[321]), .S(n26212), .Y(n28803) );
  MUX2X1 U19117 ( .B(grid[303]), .A(grid[309]), .S(n26182), .Y(n28807) );
  MUX2X1 U19118 ( .B(grid[291]), .A(grid[297]), .S(n26216), .Y(n28806) );
  MUX2X1 U19119 ( .B(n28805), .A(n28802), .S(n26550), .Y(n28809) );
  MUX2X1 U19120 ( .B(grid[279]), .A(grid[285]), .S(n26176), .Y(n28813) );
  MUX2X1 U19121 ( .B(grid[267]), .A(grid[273]), .S(n26262), .Y(n28812) );
  MUX2X1 U19122 ( .B(grid[255]), .A(grid[261]), .S(n26211), .Y(n28816) );
  MUX2X1 U19123 ( .B(grid[243]), .A(grid[249]), .S(n26174), .Y(n28815) );
  MUX2X1 U19124 ( .B(n28814), .A(n28811), .S(n26533), .Y(n28825) );
  MUX2X1 U19125 ( .B(grid[231]), .A(grid[237]), .S(n26183), .Y(n28819) );
  MUX2X1 U19126 ( .B(grid[219]), .A(grid[225]), .S(n26240), .Y(n28818) );
  MUX2X1 U19127 ( .B(grid[207]), .A(grid[213]), .S(n26238), .Y(n28822) );
  MUX2X1 U19128 ( .B(grid[195]), .A(grid[201]), .S(n26230), .Y(n28821) );
  MUX2X1 U19129 ( .B(n28820), .A(n28817), .S(n26552), .Y(n28824) );
  MUX2X1 U19130 ( .B(n28823), .A(n28808), .S(n28993), .Y(n28857) );
  MUX2X1 U19131 ( .B(grid[183]), .A(grid[189]), .S(n26253), .Y(n28828) );
  MUX2X1 U19132 ( .B(grid[171]), .A(grid[177]), .S(n26214), .Y(n28827) );
  MUX2X1 U19133 ( .B(grid[159]), .A(grid[165]), .S(n26261), .Y(n28831) );
  MUX2X1 U19134 ( .B(grid[147]), .A(grid[153]), .S(n26242), .Y(n28830) );
  MUX2X1 U19135 ( .B(n28829), .A(n28826), .S(n26549), .Y(n28840) );
  MUX2X1 U19136 ( .B(grid[135]), .A(grid[141]), .S(n26211), .Y(n28834) );
  MUX2X1 U19137 ( .B(grid[123]), .A(grid[129]), .S(n26200), .Y(n28833) );
  MUX2X1 U19138 ( .B(grid[111]), .A(grid[117]), .S(n26241), .Y(n28837) );
  MUX2X1 U19139 ( .B(grid[99]), .A(grid[105]), .S(n26202), .Y(n28836) );
  MUX2X1 U19140 ( .B(n28835), .A(n28832), .S(n26526), .Y(n28839) );
  MUX2X1 U19141 ( .B(grid[87]), .A(grid[93]), .S(n26188), .Y(n28843) );
  MUX2X1 U19142 ( .B(grid[75]), .A(grid[81]), .S(n26238), .Y(n28842) );
  MUX2X1 U19143 ( .B(grid[63]), .A(grid[69]), .S(n26241), .Y(n28846) );
  MUX2X1 U19144 ( .B(grid[51]), .A(grid[57]), .S(n26197), .Y(n28845) );
  MUX2X1 U19145 ( .B(n28844), .A(n28841), .S(n26554), .Y(n28855) );
  MUX2X1 U19146 ( .B(grid[39]), .A(grid[45]), .S(n26239), .Y(n28849) );
  MUX2X1 U19147 ( .B(grid[27]), .A(grid[33]), .S(n26201), .Y(n28848) );
  MUX2X1 U19148 ( .B(grid[15]), .A(grid[21]), .S(n26229), .Y(n28852) );
  MUX2X1 U19149 ( .B(grid[3]), .A(grid[9]), .S(n26210), .Y(n28851) );
  MUX2X1 U19150 ( .B(n28850), .A(n28847), .S(n26531), .Y(n28854) );
  MUX2X1 U19151 ( .B(n28853), .A(n28838), .S(n28993), .Y(n28856) );
  MUX2X1 U19152 ( .B(grid[376]), .A(grid[382]), .S(n26243), .Y(n28860) );
  MUX2X1 U19153 ( .B(grid[364]), .A(grid[370]), .S(n26257), .Y(n28859) );
  MUX2X1 U19154 ( .B(grid[352]), .A(grid[358]), .S(n26182), .Y(n28863) );
  MUX2X1 U19155 ( .B(grid[340]), .A(grid[346]), .S(n26227), .Y(n28862) );
  MUX2X1 U19156 ( .B(n28861), .A(n28858), .S(n26572), .Y(n28872) );
  MUX2X1 U19157 ( .B(grid[328]), .A(grid[334]), .S(n26254), .Y(n28866) );
  MUX2X1 U19158 ( .B(grid[316]), .A(grid[322]), .S(n26252), .Y(n28865) );
  MUX2X1 U19159 ( .B(grid[304]), .A(grid[310]), .S(n26225), .Y(n28869) );
  MUX2X1 U19160 ( .B(grid[292]), .A(grid[298]), .S(n26186), .Y(n28868) );
  MUX2X1 U19161 ( .B(n28867), .A(n28864), .S(n26565), .Y(n28871) );
  MUX2X1 U19162 ( .B(grid[280]), .A(grid[286]), .S(n26183), .Y(n28875) );
  MUX2X1 U19163 ( .B(grid[268]), .A(grid[274]), .S(n26228), .Y(n28874) );
  MUX2X1 U19164 ( .B(grid[256]), .A(grid[262]), .S(n26261), .Y(n28878) );
  MUX2X1 U19165 ( .B(grid[244]), .A(grid[250]), .S(n26213), .Y(n28877) );
  MUX2X1 U19166 ( .B(n28876), .A(n28873), .S(n26564), .Y(n28887) );
  MUX2X1 U19167 ( .B(grid[232]), .A(grid[238]), .S(n26265), .Y(n28881) );
  MUX2X1 U19168 ( .B(grid[220]), .A(grid[226]), .S(n26187), .Y(n28880) );
  MUX2X1 U19169 ( .B(grid[208]), .A(grid[214]), .S(n26210), .Y(n28884) );
  MUX2X1 U19170 ( .B(grid[196]), .A(grid[202]), .S(n26240), .Y(n28883) );
  MUX2X1 U19171 ( .B(n28882), .A(n28879), .S(n26566), .Y(n28886) );
  MUX2X1 U19172 ( .B(n28885), .A(n28870), .S(n28994), .Y(n28919) );
  MUX2X1 U19173 ( .B(grid[184]), .A(grid[190]), .S(n26256), .Y(n28890) );
  MUX2X1 U19174 ( .B(grid[172]), .A(grid[178]), .S(n26255), .Y(n28889) );
  MUX2X1 U19175 ( .B(grid[160]), .A(grid[166]), .S(n26177), .Y(n28893) );
  MUX2X1 U19176 ( .B(grid[148]), .A(grid[154]), .S(n26263), .Y(n28892) );
  MUX2X1 U19177 ( .B(n28891), .A(n28888), .S(n26575), .Y(n28902) );
  MUX2X1 U19178 ( .B(grid[136]), .A(grid[142]), .S(n26244), .Y(n28896) );
  MUX2X1 U19179 ( .B(grid[124]), .A(grid[130]), .S(n26213), .Y(n28895) );
  MUX2X1 U19180 ( .B(grid[112]), .A(grid[118]), .S(n26185), .Y(n28899) );
  MUX2X1 U19181 ( .B(grid[100]), .A(grid[106]), .S(n26216), .Y(n28898) );
  MUX2X1 U19182 ( .B(n28897), .A(n28894), .S(n26551), .Y(n28901) );
  MUX2X1 U19183 ( .B(grid[88]), .A(grid[94]), .S(n26226), .Y(n28905) );
  MUX2X1 U19184 ( .B(grid[76]), .A(grid[82]), .S(n26264), .Y(n28904) );
  MUX2X1 U19185 ( .B(grid[64]), .A(grid[70]), .S(n26212), .Y(n28908) );
  MUX2X1 U19186 ( .B(grid[52]), .A(grid[58]), .S(n26242), .Y(n28907) );
  MUX2X1 U19187 ( .B(n28906), .A(n28903), .S(n26574), .Y(n28917) );
  MUX2X1 U19188 ( .B(grid[40]), .A(grid[46]), .S(n26184), .Y(n28911) );
  MUX2X1 U19189 ( .B(grid[28]), .A(grid[34]), .S(n26215), .Y(n28910) );
  MUX2X1 U19190 ( .B(grid[16]), .A(grid[22]), .S(n26239), .Y(n28914) );
  MUX2X1 U19191 ( .B(grid[4]), .A(grid[10]), .S(n26196), .Y(n28913) );
  MUX2X1 U19192 ( .B(n28912), .A(n28909), .S(n26556), .Y(n28916) );
  MUX2X1 U19193 ( .B(n28915), .A(n28900), .S(n28994), .Y(n28918) );
  MUX2X1 U19194 ( .B(grid[377]), .A(grid[383]), .S(n26172), .Y(n28922) );
  MUX2X1 U19195 ( .B(grid[365]), .A(grid[371]), .S(n26187), .Y(n28921) );
  MUX2X1 U19196 ( .B(grid[353]), .A(grid[359]), .S(n26173), .Y(n28925) );
  MUX2X1 U19197 ( .B(grid[341]), .A(grid[347]), .S(n26262), .Y(n28924) );
  MUX2X1 U19198 ( .B(n28923), .A(n28920), .S(n26532), .Y(n28934) );
  MUX2X1 U19199 ( .B(grid[329]), .A(grid[335]), .S(n26186), .Y(n28928) );
  MUX2X1 U19200 ( .B(grid[317]), .A(grid[323]), .S(n26240), .Y(n28927) );
  MUX2X1 U19201 ( .B(grid[305]), .A(grid[311]), .S(n26261), .Y(n28931) );
  MUX2X1 U19202 ( .B(grid[293]), .A(grid[299]), .S(n26253), .Y(n28930) );
  MUX2X1 U19203 ( .B(n28929), .A(n28926), .S(n26539), .Y(n28933) );
  MUX2X1 U19204 ( .B(grid[281]), .A(grid[287]), .S(n26227), .Y(n28937) );
  MUX2X1 U19205 ( .B(grid[269]), .A(grid[275]), .S(n26263), .Y(n28936) );
  MUX2X1 U19206 ( .B(grid[257]), .A(grid[263]), .S(n26228), .Y(n28940) );
  MUX2X1 U19207 ( .B(grid[245]), .A(grid[251]), .S(n26267), .Y(n28939) );
  MUX2X1 U19208 ( .B(n28938), .A(n28935), .S(n26557), .Y(n28949) );
  MUX2X1 U19209 ( .B(grid[233]), .A(grid[239]), .S(n26268), .Y(n28943) );
  MUX2X1 U19210 ( .B(grid[221]), .A(grid[227]), .S(n26254), .Y(n28942) );
  MUX2X1 U19211 ( .B(grid[209]), .A(grid[215]), .S(n26266), .Y(n28946) );
  MUX2X1 U19212 ( .B(grid[197]), .A(grid[203]), .S(n26261), .Y(n28945) );
  MUX2X1 U19213 ( .B(n28944), .A(n28941), .S(n26542), .Y(n28948) );
  MUX2X1 U19214 ( .B(n28947), .A(n28932), .S(n28994), .Y(n28981) );
  MUX2X1 U19215 ( .B(grid[185]), .A(grid[191]), .S(n26188), .Y(n28952) );
  MUX2X1 U19216 ( .B(grid[173]), .A(grid[179]), .S(n26241), .Y(n28951) );
  MUX2X1 U19217 ( .B(grid[161]), .A(grid[167]), .S(n26264), .Y(n28955) );
  MUX2X1 U19218 ( .B(grid[149]), .A(grid[155]), .S(n26255), .Y(n28954) );
  MUX2X1 U19219 ( .B(n28953), .A(n28950), .S(n26538), .Y(n28964) );
  MUX2X1 U19220 ( .B(grid[137]), .A(grid[143]), .S(n26242), .Y(n28958) );
  MUX2X1 U19221 ( .B(grid[125]), .A(grid[131]), .S(n26253), .Y(n28957) );
  MUX2X1 U19222 ( .B(grid[113]), .A(grid[119]), .S(n26256), .Y(n28961) );
  MUX2X1 U19223 ( .B(grid[101]), .A(grid[107]), .S(n26263), .Y(n28960) );
  MUX2X1 U19224 ( .B(n28959), .A(n28956), .S(n26537), .Y(n28963) );
  MUX2X1 U19225 ( .B(grid[89]), .A(grid[95]), .S(n26265), .Y(n28967) );
  MUX2X1 U19226 ( .B(grid[77]), .A(grid[83]), .S(n26258), .Y(n28966) );
  MUX2X1 U19227 ( .B(grid[65]), .A(grid[71]), .S(n26268), .Y(n28970) );
  MUX2X1 U19228 ( .B(grid[53]), .A(grid[59]), .S(n26262), .Y(n28969) );
  MUX2X1 U19229 ( .B(n28968), .A(n28965), .S(n26541), .Y(n28979) );
  MUX2X1 U19230 ( .B(grid[41]), .A(grid[47]), .S(n26257), .Y(n28973) );
  MUX2X1 U19231 ( .B(grid[29]), .A(grid[35]), .S(n26264), .Y(n28972) );
  MUX2X1 U19232 ( .B(grid[17]), .A(grid[23]), .S(n26184), .Y(n28976) );
  MUX2X1 U19233 ( .B(grid[5]), .A(grid[11]), .S(n26202), .Y(n28975) );
  MUX2X1 U19234 ( .B(n28974), .A(n28971), .S(n26540), .Y(n28978) );
  MUX2X1 U19235 ( .B(n28977), .A(n28962), .S(n28994), .Y(n28980) );
  MUX2X1 U19236 ( .B(n28996), .A(n28997), .S(n29182), .Y(n28995) );
  MUX2X1 U19237 ( .B(n28999), .A(n29000), .S(n29182), .Y(n28998) );
  MUX2X1 U19238 ( .B(n29002), .A(n29003), .S(n29182), .Y(n29001) );
  MUX2X1 U19239 ( .B(n29005), .A(n29006), .S(n29182), .Y(n29004) );
  MUX2X1 U19240 ( .B(n29008), .A(n29009), .S(n29186), .Y(n29007) );
  MUX2X1 U19241 ( .B(n29011), .A(n29012), .S(n29181), .Y(n29010) );
  MUX2X1 U19242 ( .B(n29014), .A(n29015), .S(n29182), .Y(n29013) );
  MUX2X1 U19243 ( .B(n29017), .A(n29018), .S(n29182), .Y(n29016) );
  MUX2X1 U19244 ( .B(n29020), .A(n29021), .S(n29182), .Y(n29019) );
  MUX2X1 U19245 ( .B(n29023), .A(n29024), .S(n29187), .Y(n29022) );
  MUX2X1 U19246 ( .B(n29026), .A(n29027), .S(n29182), .Y(n29025) );
  MUX2X1 U19247 ( .B(n29029), .A(n29030), .S(n29182), .Y(n29028) );
  MUX2X1 U19248 ( .B(n29032), .A(n29033), .S(n29182), .Y(n29031) );
  MUX2X1 U19249 ( .B(n29035), .A(n29036), .S(n29182), .Y(n29034) );
  MUX2X1 U19250 ( .B(n29038), .A(n29039), .S(n29186), .Y(n29037) );
  MUX2X1 U19251 ( .B(n29041), .A(n29042), .S(n29182), .Y(n29040) );
  MUX2X1 U19252 ( .B(n29044), .A(n29045), .S(n29182), .Y(n29043) );
  MUX2X1 U19253 ( .B(n29047), .A(n29048), .S(n29182), .Y(n29046) );
  MUX2X1 U19254 ( .B(n29050), .A(n29051), .S(n29182), .Y(n29049) );
  MUX2X1 U19255 ( .B(n29053), .A(n29054), .S(n29187), .Y(n29052) );
  MUX2X1 U19256 ( .B(n25472), .A(n29055), .S(n2256), .Y(n19664) );
  MUX2X1 U19257 ( .B(n29057), .A(n29058), .S(n29182), .Y(n29056) );
  MUX2X1 U19258 ( .B(n29060), .A(n29061), .S(n29182), .Y(n29059) );
  MUX2X1 U19259 ( .B(n29063), .A(n29064), .S(n29182), .Y(n29062) );
  MUX2X1 U19260 ( .B(n29066), .A(n29067), .S(n29182), .Y(n29065) );
  MUX2X1 U19261 ( .B(n29069), .A(n29070), .S(n29186), .Y(n29068) );
  MUX2X1 U19262 ( .B(n29072), .A(n29073), .S(n29182), .Y(n29071) );
  MUX2X1 U19263 ( .B(n29075), .A(n29076), .S(n29181), .Y(n29074) );
  MUX2X1 U19264 ( .B(n29078), .A(n29079), .S(n29182), .Y(n29077) );
  MUX2X1 U19265 ( .B(n29081), .A(n29082), .S(n29182), .Y(n29080) );
  MUX2X1 U19266 ( .B(n29084), .A(n25527), .S(n29187), .Y(n29083) );
  MUX2X1 U19267 ( .B(n29086), .A(n29087), .S(n29182), .Y(n29085) );
  MUX2X1 U19268 ( .B(n29089), .A(n29090), .S(n29182), .Y(n29088) );
  MUX2X1 U19269 ( .B(n29092), .A(n29093), .S(n29182), .Y(n29091) );
  MUX2X1 U19270 ( .B(n29095), .A(n29096), .S(n29182), .Y(n29094) );
  MUX2X1 U19271 ( .B(n29098), .A(n29099), .S(n29186), .Y(n29097) );
  MUX2X1 U19272 ( .B(n29101), .A(n29102), .S(n29182), .Y(n29100) );
  MUX2X1 U19273 ( .B(n29104), .A(n29105), .S(n29182), .Y(n29103) );
  MUX2X1 U19274 ( .B(n29107), .A(n29108), .S(n29182), .Y(n29106) );
  MUX2X1 U19275 ( .B(n29110), .A(n29111), .S(n29182), .Y(n29109) );
  MUX2X1 U19276 ( .B(n29113), .A(n29114), .S(n29187), .Y(n29112) );
  MUX2X1 U19277 ( .B(n29115), .A(n25524), .S(n2256), .Y(n19663) );
  MUX2X1 U19278 ( .B(n29117), .A(n29118), .S(n29181), .Y(n29116) );
  MUX2X1 U19279 ( .B(n29120), .A(n29121), .S(n29180), .Y(n29119) );
  MUX2X1 U19280 ( .B(n29123), .A(n29124), .S(n29181), .Y(n29122) );
  MUX2X1 U19281 ( .B(n29126), .A(n29127), .S(n29181), .Y(n29125) );
  MUX2X1 U19282 ( .B(n29129), .A(n29130), .S(n29186), .Y(n29128) );
  MUX2X1 U19283 ( .B(n29132), .A(n29133), .S(n29182), .Y(n29131) );
  MUX2X1 U19284 ( .B(n29135), .A(n29136), .S(n29182), .Y(n29134) );
  MUX2X1 U19285 ( .B(n29138), .A(n29139), .S(n29182), .Y(n29137) );
  MUX2X1 U19286 ( .B(n29141), .A(n29142), .S(n29182), .Y(n29140) );
  MUX2X1 U19287 ( .B(n29144), .A(n29145), .S(n29187), .Y(n29143) );
  MUX2X1 U19288 ( .B(n29147), .A(n29148), .S(n29180), .Y(n29146) );
  MUX2X1 U19289 ( .B(n29150), .A(n29151), .S(n29181), .Y(n29149) );
  MUX2X1 U19290 ( .B(n29153), .A(n29154), .S(n29182), .Y(n29152) );
  MUX2X1 U19291 ( .B(n29156), .A(n29157), .S(n29182), .Y(n29155) );
  MUX2X1 U19292 ( .B(n29159), .A(n29160), .S(n29186), .Y(n29158) );
  MUX2X1 U19293 ( .B(n29162), .A(n29163), .S(n29180), .Y(n29161) );
  MUX2X1 U19294 ( .B(n29168), .A(n29169), .S(n29181), .Y(n29167) );
  MUX2X1 U19295 ( .B(n29171), .A(n29172), .S(n29180), .Y(n29170) );
  MUX2X1 U19296 ( .B(n29174), .A(n29175), .S(n29187), .Y(n29173) );
  MUX2X1 U19297 ( .B(n29176), .A(n29177), .S(n2256), .Y(n19662) );
  MUX2X1 U19298 ( .B(grid[372]), .A(grid[378]), .S(net150650), .Y(n28997) );
  MUX2X1 U19299 ( .B(grid[360]), .A(grid[366]), .S(alt5_net95664), .Y(n28996)
         );
  MUX2X1 U19300 ( .B(grid[348]), .A(grid[354]), .S(net150650), .Y(n29000) );
  MUX2X1 U19301 ( .B(grid[336]), .A(grid[342]), .S(net150650), .Y(n28999) );
  MUX2X1 U19302 ( .B(n28998), .A(n28995), .S(n29185), .Y(n29009) );
  MUX2X1 U19303 ( .B(grid[324]), .A(grid[330]), .S(alt5_net95652), .Y(n29003)
         );
  MUX2X1 U19304 ( .B(grid[312]), .A(grid[318]), .S(net113321), .Y(n29002) );
  MUX2X1 U19305 ( .B(grid[300]), .A(grid[306]), .S(net113321), .Y(n29006) );
  MUX2X1 U19306 ( .B(grid[288]), .A(grid[294]), .S(alt5_net95652), .Y(n29005)
         );
  MUX2X1 U19307 ( .B(n29004), .A(n29001), .S(n29185), .Y(n29008) );
  MUX2X1 U19308 ( .B(grid[276]), .A(grid[282]), .S(alt5_net95664), .Y(n29012)
         );
  MUX2X1 U19309 ( .B(grid[264]), .A(grid[270]), .S(alt5_net95666), .Y(n29011)
         );
  MUX2X1 U19310 ( .B(grid[252]), .A(grid[258]), .S(alt5_net95664), .Y(n29015)
         );
  MUX2X1 U19311 ( .B(grid[240]), .A(grid[246]), .S(alt5_net95664), .Y(n29014)
         );
  MUX2X1 U19312 ( .B(n29013), .A(n29010), .S(n29185), .Y(n29024) );
  MUX2X1 U19313 ( .B(grid[228]), .A(grid[234]), .S(alt5_net95654), .Y(n29018)
         );
  MUX2X1 U19314 ( .B(grid[216]), .A(grid[222]), .S(alt5_net95654), .Y(n29017)
         );
  MUX2X1 U19315 ( .B(grid[204]), .A(grid[210]), .S(alt5_net95654), .Y(n29021)
         );
  MUX2X1 U19316 ( .B(grid[192]), .A(grid[198]), .S(alt5_net95654), .Y(n29020)
         );
  MUX2X1 U19317 ( .B(n29019), .A(n29016), .S(n29185), .Y(n29023) );
  MUX2X1 U19318 ( .B(n29022), .A(n29007), .S(n2255), .Y(n29055) );
  MUX2X1 U19319 ( .B(grid[180]), .A(grid[186]), .S(alt5_net95654), .Y(n29027)
         );
  MUX2X1 U19320 ( .B(grid[168]), .A(grid[174]), .S(alt5_net95654), .Y(n29026)
         );
  MUX2X1 U19321 ( .B(grid[156]), .A(grid[162]), .S(alt5_net95654), .Y(n29030)
         );
  MUX2X1 U19322 ( .B(grid[144]), .A(grid[150]), .S(alt5_net95654), .Y(n29029)
         );
  MUX2X1 U19323 ( .B(n29028), .A(n29025), .S(n29185), .Y(n29039) );
  MUX2X1 U19324 ( .B(grid[132]), .A(grid[138]), .S(alt5_net95654), .Y(n29033)
         );
  MUX2X1 U19325 ( .B(grid[120]), .A(grid[126]), .S(alt5_net95654), .Y(n29032)
         );
  MUX2X1 U19326 ( .B(grid[108]), .A(grid[114]), .S(alt5_net95654), .Y(n29036)
         );
  MUX2X1 U19327 ( .B(grid[96]), .A(grid[102]), .S(alt5_net95654), .Y(n29035)
         );
  MUX2X1 U19328 ( .B(n29034), .A(n29031), .S(n29185), .Y(n29038) );
  MUX2X1 U19329 ( .B(grid[84]), .A(grid[90]), .S(alt5_net95656), .Y(n29042) );
  MUX2X1 U19330 ( .B(grid[72]), .A(grid[78]), .S(alt5_net95656), .Y(n29041) );
  MUX2X1 U19331 ( .B(grid[60]), .A(grid[66]), .S(alt5_net95656), .Y(n29045) );
  MUX2X1 U19332 ( .B(grid[48]), .A(grid[54]), .S(alt5_net95656), .Y(n29044) );
  MUX2X1 U19333 ( .B(n29043), .A(n29040), .S(n29185), .Y(n29054) );
  MUX2X1 U19334 ( .B(grid[36]), .A(grid[42]), .S(alt5_net95656), .Y(n29048) );
  MUX2X1 U19335 ( .B(grid[24]), .A(grid[30]), .S(alt5_net95656), .Y(n29047) );
  MUX2X1 U19336 ( .B(grid[12]), .A(grid[18]), .S(alt5_net95656), .Y(n29051) );
  MUX2X1 U19337 ( .B(grid[0]), .A(grid[6]), .S(alt5_net95656), .Y(n29050) );
  MUX2X1 U19338 ( .B(n29049), .A(n29046), .S(n29185), .Y(n29053) );
  MUX2X1 U19339 ( .B(grid[373]), .A(grid[379]), .S(alt5_net95656), .Y(n29058)
         );
  MUX2X1 U19340 ( .B(grid[361]), .A(grid[367]), .S(alt5_net95656), .Y(n29057)
         );
  MUX2X1 U19341 ( .B(grid[349]), .A(grid[355]), .S(alt5_net95656), .Y(n29061)
         );
  MUX2X1 U19342 ( .B(grid[337]), .A(grid[343]), .S(alt5_net95656), .Y(n29060)
         );
  MUX2X1 U19343 ( .B(n29059), .A(n29056), .S(n29185), .Y(n29070) );
  MUX2X1 U19344 ( .B(grid[325]), .A(grid[331]), .S(alt5_net95658), .Y(n29064)
         );
  MUX2X1 U19345 ( .B(grid[313]), .A(grid[319]), .S(alt5_net95658), .Y(n29063)
         );
  MUX2X1 U19346 ( .B(grid[301]), .A(grid[307]), .S(alt5_net95658), .Y(n29067)
         );
  MUX2X1 U19347 ( .B(grid[289]), .A(grid[295]), .S(alt5_net95658), .Y(n29066)
         );
  MUX2X1 U19348 ( .B(n29065), .A(n29062), .S(n29185), .Y(n29069) );
  MUX2X1 U19349 ( .B(grid[277]), .A(grid[283]), .S(alt5_net95658), .Y(n29073)
         );
  MUX2X1 U19350 ( .B(grid[265]), .A(grid[271]), .S(alt5_net95658), .Y(n29072)
         );
  MUX2X1 U19351 ( .B(grid[253]), .A(grid[259]), .S(alt5_net95658), .Y(n29076)
         );
  MUX2X1 U19352 ( .B(grid[241]), .A(grid[247]), .S(alt5_net95658), .Y(n29075)
         );
  MUX2X1 U19353 ( .B(grid[229]), .A(grid[235]), .S(alt5_net95658), .Y(n29079)
         );
  MUX2X1 U19354 ( .B(grid[217]), .A(grid[223]), .S(alt5_net95658), .Y(n29078)
         );
  MUX2X1 U19355 ( .B(grid[205]), .A(grid[211]), .S(alt5_net95658), .Y(n29082)
         );
  MUX2X1 U19356 ( .B(grid[193]), .A(grid[199]), .S(alt5_net95658), .Y(n29081)
         );
  MUX2X1 U19357 ( .B(n29080), .A(n29077), .S(n29185), .Y(n29084) );
  MUX2X1 U19358 ( .B(grid[181]), .A(grid[187]), .S(alt5_net95662), .Y(n29087)
         );
  MUX2X1 U19359 ( .B(grid[169]), .A(grid[175]), .S(net150650), .Y(n29086) );
  MUX2X1 U19360 ( .B(grid[157]), .A(grid[163]), .S(alt5_net95666), .Y(n29090)
         );
  MUX2X1 U19361 ( .B(grid[145]), .A(grid[151]), .S(alt5_net95662), .Y(n29089)
         );
  MUX2X1 U19362 ( .B(n29088), .A(n29085), .S(n29184), .Y(n29099) );
  MUX2X1 U19363 ( .B(grid[133]), .A(grid[139]), .S(alt5_net95666), .Y(n29093)
         );
  MUX2X1 U19364 ( .B(grid[121]), .A(grid[127]), .S(net150650), .Y(n29092) );
  MUX2X1 U19365 ( .B(grid[109]), .A(grid[115]), .S(net113321), .Y(n29096) );
  MUX2X1 U19366 ( .B(grid[97]), .A(grid[103]), .S(alt5_net95652), .Y(n29095)
         );
  MUX2X1 U19367 ( .B(n29094), .A(n29091), .S(n29184), .Y(n29098) );
  MUX2X1 U19368 ( .B(grid[85]), .A(grid[91]), .S(net150650), .Y(n29102) );
  MUX2X1 U19369 ( .B(grid[73]), .A(grid[79]), .S(alt5_net95666), .Y(n29101) );
  MUX2X1 U19370 ( .B(grid[61]), .A(grid[67]), .S(alt5_net95662), .Y(n29105) );
  MUX2X1 U19371 ( .B(grid[49]), .A(grid[55]), .S(net150650), .Y(n29104) );
  MUX2X1 U19372 ( .B(n29103), .A(n29100), .S(n29184), .Y(n29114) );
  MUX2X1 U19373 ( .B(grid[37]), .A(grid[43]), .S(alt5_net95664), .Y(n29108) );
  MUX2X1 U19374 ( .B(grid[25]), .A(grid[31]), .S(net150650), .Y(n29107) );
  MUX2X1 U19375 ( .B(grid[13]), .A(grid[19]), .S(alt5_net95662), .Y(n29111) );
  MUX2X1 U19376 ( .B(grid[1]), .A(grid[7]), .S(alt5_net95666), .Y(n29110) );
  MUX2X1 U19377 ( .B(n29109), .A(n29106), .S(n29184), .Y(n29113) );
  MUX2X1 U19378 ( .B(n29112), .A(n29097), .S(n2255), .Y(n29115) );
  MUX2X1 U19379 ( .B(grid[374]), .A(grid[380]), .S(net150650), .Y(n29118) );
  MUX2X1 U19380 ( .B(grid[362]), .A(grid[368]), .S(net150650), .Y(n29117) );
  MUX2X1 U19381 ( .B(grid[350]), .A(grid[356]), .S(net150650), .Y(n29121) );
  MUX2X1 U19382 ( .B(grid[338]), .A(grid[344]), .S(alt5_net95666), .Y(n29120)
         );
  MUX2X1 U19383 ( .B(n29119), .A(n29116), .S(n29184), .Y(n29130) );
  MUX2X1 U19384 ( .B(grid[326]), .A(grid[332]), .S(alt5_net95666), .Y(n29124)
         );
  MUX2X1 U19385 ( .B(grid[314]), .A(grid[320]), .S(alt5_net95664), .Y(n29123)
         );
  MUX2X1 U19386 ( .B(grid[302]), .A(grid[308]), .S(net150650), .Y(n29127) );
  MUX2X1 U19387 ( .B(grid[290]), .A(grid[296]), .S(alt5_net95662), .Y(n29126)
         );
  MUX2X1 U19388 ( .B(n29125), .A(n29122), .S(n29184), .Y(n29129) );
  MUX2X1 U19389 ( .B(grid[278]), .A(grid[284]), .S(net113321), .Y(n29133) );
  MUX2X1 U19390 ( .B(grid[266]), .A(grid[272]), .S(alt5_net95666), .Y(n29132)
         );
  MUX2X1 U19391 ( .B(grid[254]), .A(grid[260]), .S(alt5_net95666), .Y(n29136)
         );
  MUX2X1 U19392 ( .B(grid[242]), .A(grid[248]), .S(alt5_net95664), .Y(n29135)
         );
  MUX2X1 U19393 ( .B(n29134), .A(n29131), .S(n29184), .Y(n29145) );
  MUX2X1 U19394 ( .B(grid[230]), .A(grid[236]), .S(net150650), .Y(n29139) );
  MUX2X1 U19395 ( .B(grid[218]), .A(grid[224]), .S(net150650), .Y(n29138) );
  MUX2X1 U19396 ( .B(grid[206]), .A(grid[212]), .S(alt5_net95652), .Y(n29142)
         );
  MUX2X1 U19397 ( .B(grid[194]), .A(grid[200]), .S(alt5_net95666), .Y(n29141)
         );
  MUX2X1 U19398 ( .B(n29140), .A(n29137), .S(n29184), .Y(n29144) );
  MUX2X1 U19399 ( .B(n29143), .A(n29128), .S(n2255), .Y(n29177) );
  MUX2X1 U19400 ( .B(grid[182]), .A(grid[188]), .S(net150650), .Y(n29148) );
  MUX2X1 U19401 ( .B(grid[170]), .A(grid[176]), .S(net150650), .Y(n29147) );
  MUX2X1 U19402 ( .B(grid[158]), .A(grid[164]), .S(net113321), .Y(n29151) );
  MUX2X1 U19403 ( .B(grid[146]), .A(grid[152]), .S(alt5_net95664), .Y(n29150)
         );
  MUX2X1 U19404 ( .B(n29149), .A(n29146), .S(n29184), .Y(n29160) );
  MUX2X1 U19405 ( .B(grid[134]), .A(grid[140]), .S(alt5_net95652), .Y(n29154)
         );
  MUX2X1 U19406 ( .B(grid[122]), .A(grid[128]), .S(alt5_net95664), .Y(n29153)
         );
  MUX2X1 U19407 ( .B(grid[110]), .A(grid[116]), .S(net150650), .Y(n29157) );
  MUX2X1 U19408 ( .B(grid[98]), .A(grid[104]), .S(alt5_net95662), .Y(n29156)
         );
  MUX2X1 U19409 ( .B(n29155), .A(n29152), .S(n29184), .Y(n29159) );
  MUX2X1 U19410 ( .B(grid[86]), .A(grid[92]), .S(net150650), .Y(n29163) );
  MUX2X1 U19411 ( .B(grid[74]), .A(grid[80]), .S(alt5_net95664), .Y(n29162) );
  MUX2X1 U19412 ( .B(grid[62]), .A(grid[68]), .S(net150650), .Y(n29166) );
  MUX2X1 U19413 ( .B(grid[50]), .A(grid[56]), .S(alt5_net95652), .Y(n29165) );
  MUX2X1 U19414 ( .B(n29164), .A(n29161), .S(n29184), .Y(n29175) );
  MUX2X1 U19415 ( .B(grid[38]), .A(grid[44]), .S(net150650), .Y(n29169) );
  MUX2X1 U19416 ( .B(grid[26]), .A(grid[32]), .S(net113321), .Y(n29168) );
  MUX2X1 U19417 ( .B(grid[14]), .A(grid[20]), .S(alt5_net95664), .Y(n29172) );
  MUX2X1 U19418 ( .B(grid[2]), .A(grid[8]), .S(alt5_net95666), .Y(n29171) );
  MUX2X1 U19419 ( .B(n29170), .A(n29167), .S(n29184), .Y(n29174) );
  MUX2X1 U19420 ( .B(n29173), .A(n29158), .S(n2255), .Y(n29176) );
  INVX1 U19421 ( .A(nc[5]), .Y(n29540) );
  INVX1 U19422 ( .A(nc[13]), .Y(n29544) );
  AND2X1 U19423 ( .A(n9144), .B(n29381), .Y(n21802) );
  AND2X1 U19424 ( .A(n9142), .B(n29381), .Y(n21799) );
  AND2X1 U19425 ( .A(n9140), .B(n29381), .Y(n21797) );
  AND2X1 U19426 ( .A(n9138), .B(n29381), .Y(n21795) );
  AND2X1 U19427 ( .A(n9132), .B(n29381), .Y(n21789) );
  INVX1 U19428 ( .A(n26788), .Y(n29730) );
  INVX1 U19429 ( .A(n23067), .Y(n30637) );
  INVX1 U19430 ( .A(n23125), .Y(n31368) );
  INVX1 U19431 ( .A(n23123), .Y(n31348) );
  INVX1 U19432 ( .A(n23198), .Y(n31328) );
  INVX1 U19433 ( .A(n23167), .Y(n31254) );
  INVX1 U19434 ( .A(n23165), .Y(n31214) );
  INVX1 U19435 ( .A(n23122), .Y(n31137) );
  INVX1 U19436 ( .A(n23131), .Y(n31836) );
  INVX1 U19437 ( .A(n22980), .Y(n29513) );
  INVX1 U19438 ( .A(net125067), .Y(net95105) );
  INVX1 U19439 ( .A(n23075), .Y(n30632) );
  INVX1 U19440 ( .A(n33000), .Y(n33058) );
  INVX1 U19441 ( .A(n23080), .Y(n33057) );
  AND2X2 U19442 ( .A(n23291), .B(n21106), .Y(n29190) );
  NOR3X1 U19443 ( .A(locTrig[1]), .B(n21059), .C(n29192), .Y(n29191) );
  INVX1 U19444 ( .A(n26278), .Y(n29194) );
  INVX1 U19445 ( .A(n23138), .Y(n31468) );
  INVX1 U19446 ( .A(n22965), .Y(n29196) );
  INVX1 U19447 ( .A(n29220), .Y(n29219) );
  INVX1 U19448 ( .A(n22965), .Y(n29220) );
  INVX1 U19449 ( .A(n23121), .Y(n30962) );
  INVX1 U19450 ( .A(n23194), .Y(n30941) );
  INVX1 U19451 ( .A(n23119), .Y(n30922) );
  INVX1 U19452 ( .A(n23134), .Y(n30901) );
  INVX1 U19453 ( .A(n23077), .Y(n30881) );
  INVX1 U19454 ( .A(n31901), .Y(n29204) );
  INVX1 U19455 ( .A(n29199), .Y(n31857) );
  INVX1 U19456 ( .A(n29201), .Y(n31740) );
  INVX1 U19457 ( .A(n29202), .Y(n31626) );
  INVX1 U19458 ( .A(n29200), .Y(n31158) );
  INVX1 U19459 ( .A(n29198), .Y(n31040) );
  INVX1 U19460 ( .A(n29203), .Y(n31002) );
  AOI21X1 U19461 ( .A(n32287), .B(n29197), .C(n27231), .Y(n29198) );
  AOI21X1 U19462 ( .A(n23420), .B(n29197), .C(n27229), .Y(n29199) );
  AOI21X1 U19463 ( .A(n32311), .B(n29197), .C(n27228), .Y(n29200) );
  AOI21X1 U19464 ( .A(n23407), .B(n29197), .C(n27227), .Y(n29201) );
  AOI21X1 U19465 ( .A(n32407), .B(n29197), .C(n27226), .Y(n29202) );
  AOI21X1 U19466 ( .A(n32279), .B(n29197), .C(n27230), .Y(n29203) );
  INVX1 U19467 ( .A(n29208), .Y(n29233) );
  INVX1 U19468 ( .A(n29208), .Y(n29205) );
  INVX1 U19469 ( .A(n12058), .Y(n33267) );
  INVX1 U19470 ( .A(n12030), .Y(n33412) );
  INVX1 U19471 ( .A(n12036), .Y(n33382) );
  INVX1 U19472 ( .A(n12052), .Y(n33298) );
  INVX1 U19473 ( .A(n12054), .Y(n33290) );
  XOR2X1 U19474 ( .A(n33145), .B(n33146), .Y(n29206) );
  INVX1 U19475 ( .A(n12060), .Y(n33260) );
  INVX1 U19476 ( .A(n8035), .Y(n30047) );
  INVX1 U19477 ( .A(n32846), .Y(n33049) );
  INVX1 U19478 ( .A(n32657), .Y(n33053) );
  INVX1 U19479 ( .A(n21024), .Y(n29492) );
  INVX1 U19480 ( .A(n25078), .Y(n30064) );
  INVX1 U19481 ( .A(n34313), .Y(n33175) );
  INVX1 U19482 ( .A(n32612), .Y(n33054) );
  NAND3X1 U19483 ( .A(net108478), .B(net109385), .C(net115619), .Y(n14358) );
  NAND3X1 U19484 ( .A(net109512), .B(net108471), .C(net111332), .Y(n14357) );
  MUX2X1 U19485 ( .B(n25772), .A(net94649), .S(n27296), .Y(n29472) );
  OAI21X1 U19486 ( .A(net151887), .B(n26075), .C(n29472), .Y(net90071) );
  XOR2X1 U19487 ( .A(n24925), .B(n2253), .Y(n34187) );
  OAI21X1 U19488 ( .A(n27302), .B(n29465), .C(n27083), .Y(n34185) );
  AOI22X1 U19489 ( .A(n29185), .B(n23141), .C(n26164), .D(n25593), .Y(n29474)
         );
  OAI21X1 U19490 ( .A(net110410), .B(n34187), .C(n21561), .Y(net89777) );
  XOR2X1 U19491 ( .A(n29504), .B(n2254), .Y(net89744) );
  INVX2 U19492 ( .A(n2254), .Y(n34210) );
  AOI22X1 U19493 ( .A(n34210), .B(n23142), .C(n25731), .D(n25593), .Y(net95464) );
  OAI21X1 U19494 ( .A(net110410), .B(net89744), .C(net142478), .Y(n34215) );
  INVX2 U19495 ( .A(n2255), .Y(n29476) );
  MUX2X1 U19496 ( .B(n2255), .A(n29509), .S(n29477), .Y(n29478) );
  AOI22X1 U19497 ( .A(n27318), .B(net94649), .C(n27186), .D(n25836), .Y(
        net95456) );
  MUX2X1 U19498 ( .B(net94645), .A(net94647), .S(n27297), .Y(net95457) );
  AOI22X1 U19499 ( .A(n27321), .B(net94647), .C(n27317), .D(net110411), .Y(
        n29483) );
  OAI21X1 U19500 ( .A(n27256), .B(n29508), .C(n21191), .Y(n34197) );
  AOI22X1 U19501 ( .A(n34197), .B(n25593), .C(n27320), .D(net94645), .Y(n29482) );
  NAND3X1 U19502 ( .A(n29602), .B(n21192), .C(locTrig[0]), .Y(n30652) );
  AOI21X1 U19503 ( .A(direction_lee[1]), .B(n21125), .C(n24980), .Y(n29485) );
  NAND3X1 U19504 ( .A(n29490), .B(n21013), .C(n21031), .Y(n15186) );
  NAND3X1 U19505 ( .A(n21024), .B(n21101), .C(n29491), .Y(n15184) );
  NAND3X1 U19506 ( .A(n29492), .B(n21101), .C(n21028), .Y(n15179) );
  MUX2X1 U19507 ( .B(n29507), .A(n29506), .S(n27296), .Y(n29494) );
  OAI21X1 U19508 ( .A(n21074), .B(n26076), .C(n29494), .Y(n8051) );
  AOI22X1 U19509 ( .A(n29185), .B(n29496), .C(n26164), .D(n23465), .Y(n29495)
         );
  OAI21X1 U19510 ( .A(n25663), .B(n34187), .C(n21562), .Y(n8052) );
  AOI22X1 U19511 ( .A(n25777), .B(n34210), .C(n25731), .D(n23465), .Y(n29497)
         );
  OAI21X1 U19512 ( .A(n25663), .B(net89744), .C(n21563), .Y(n8053) );
  AOI22X1 U19513 ( .A(n27318), .B(n29506), .C(n27186), .D(n23465), .Y(n29499)
         );
  MUX2X1 U19514 ( .B(n29513), .A(n29511), .S(n27297), .Y(n29498) );
  AOI22X1 U19515 ( .A(n27321), .B(n29511), .C(n27317), .D(n29506), .Y(n29501)
         );
  AOI22X1 U19516 ( .A(n34197), .B(n23465), .C(n27320), .D(n29513), .Y(n29500)
         );
  NOR3X1 U19517 ( .A(n22933), .B(n21194), .C(n29508), .Y(n29517) );
  AOI21X1 U19518 ( .A(n24266), .B(n23465), .C(n29506), .Y(n29516) );
  AOI22X1 U19519 ( .A(n24328), .B(n29513), .C(n24695), .D(n29511), .Y(n29515)
         );
  OAI21X1 U19520 ( .A(n29517), .B(n24684), .C(n23748), .Y(n30066) );
  XOR2X1 U19521 ( .A(S[1]), .B(n29181), .Y(n29520) );
  XOR2X1 U19522 ( .A(S[4]), .B(n2255), .Y(n29519) );
  XOR2X1 U19523 ( .A(S[5]), .B(n2256), .Y(n29518) );
  NOR3X1 U19524 ( .A(n29520), .B(n29519), .C(n29518), .Y(n29525) );
  XOR2X1 U19525 ( .A(S[2]), .B(n29185), .Y(n29523) );
  XOR2X1 U19526 ( .A(S[0]), .B(net150650), .Y(n29522) );
  XOR2X1 U19527 ( .A(S[3]), .B(n2254), .Y(n29521) );
  NOR3X1 U19528 ( .A(n29523), .B(n29522), .C(n29521), .Y(n29524) );
  NOR3X1 U19529 ( .A(nc[28]), .B(nc[29]), .C(nc[30]), .Y(n29539) );
  NAND3X1 U19530 ( .A(n29530), .B(n26901), .C(n29528), .Y(n29535) );
  NAND3X1 U19531 ( .A(n29533), .B(n26667), .C(n29531), .Y(n29534) );
  NOR3X1 U19532 ( .A(nc[24]), .B(nc[25]), .C(n29536), .Y(n29537) );
  NAND3X1 U19533 ( .A(n29539), .B(n22728), .C(n29537), .Y(n29556) );
  NAND3X1 U19534 ( .A(n29542), .B(n26840), .C(n29540), .Y(n29548) );
  NOR3X1 U19535 ( .A(nc[14]), .B(nc[0]), .C(nc[15]), .Y(n29545) );
  NAND3X1 U19536 ( .A(n29545), .B(n29544), .C(n26737), .Y(n29546) );
  NOR3X1 U19537 ( .A(n26839), .B(n29547), .C(n26736), .Y(n29553) );
  AOI21X1 U19538 ( .A(n29553), .B(n21366), .C(nc[31]), .Y(n29554) );
  AOI21X1 U19539 ( .A(n24256), .B(n29555), .C(n22145), .Y(n29557) );
  NAND3X1 U19540 ( .A(direct[2]), .B(n29558), .C(n29559), .Y(n30650) );
  NAND3X1 U19541 ( .A(direct[1]), .B(n29560), .C(n29558), .Y(n29583) );
  NAND3X1 U19542 ( .A(direct[0]), .B(n29560), .C(n29559), .Y(n30651) );
  NAND3X1 U19543 ( .A(direct[0]), .B(direct[1]), .C(n29560), .Y(n30633) );
  MUX2X1 U19544 ( .B(n27300), .A(n29565), .S(n20813), .Y(n13703) );
  AOI21X1 U19545 ( .A(loc_s2[0]), .B(n33993), .C(n13703), .Y(n29561) );
  MUX2X1 U19546 ( .B(n29565), .A(n27300), .S(n30127), .Y(n2245) );
  OAI21X1 U19547 ( .A(n29565), .B(n26074), .C(n29562), .Y(n13704) );
  AOI21X1 U19548 ( .A(loc_s2[1]), .B(n33993), .C(n13704), .Y(n29563) );
  MUX2X1 U19549 ( .B(n34503), .A(n29595), .S(n30127), .Y(n29564) );
  MUX2X1 U19550 ( .B(n23143), .A(n21369), .S(n29683), .Y(n29567) );
  OAI21X1 U19551 ( .A(n29207), .B(n27160), .C(n29567), .Y(n2246) );
  AOI22X1 U19552 ( .A(n2253), .B(n25409), .C(n34503), .D(n34185), .Y(n29568)
         );
  OAI21X1 U19553 ( .A(n29207), .B(n34187), .C(n21564), .Y(n13705) );
  AOI21X1 U19554 ( .A(loc_s2[2]), .B(n33993), .C(n13705), .Y(n29569) );
  MUX2X1 U19555 ( .B(n27196), .A(n29207), .S(n29683), .Y(n29571) );
  OAI21X1 U19556 ( .A(n29571), .B(n23144), .C(n23441), .Y(n29573) );
  NAND3X1 U19557 ( .A(n34189), .B(n23611), .C(n21007), .Y(n29662) );
  NAND3X1 U19558 ( .A(n23102), .B(n29573), .C(n24868), .Y(n2247) );
  AOI22X1 U19559 ( .A(n25409), .B(n34210), .C(n27319), .D(n34503), .Y(n29574)
         );
  OAI21X1 U19560 ( .A(n29207), .B(net89744), .C(n21565), .Y(n13706) );
  XOR2X1 U19561 ( .A(n27176), .B(n21184), .Y(n29676) );
  AOI22X1 U19562 ( .A(n20977), .B(n25409), .C(n34503), .D(n29676), .Y(n29576)
         );
  OAI21X1 U19563 ( .A(n27254), .B(n29207), .C(n21566), .Y(n2248) );
  AOI22X1 U19564 ( .A(n27318), .B(n29595), .C(n34503), .D(n27186), .Y(n29578)
         );
  MUX2X1 U19565 ( .B(n29628), .A(n29629), .S(n27297), .Y(n29577) );
  MUX2X1 U19566 ( .B(n29590), .A(n29579), .S(n21184), .Y(n29580) );
  OAI21X1 U19567 ( .A(n26163), .B(n27196), .C(n21143), .Y(n29582) );
  OAI21X1 U19568 ( .A(n29207), .B(n25420), .C(n25335), .Y(n29586) );
  MUX2X1 U19569 ( .B(n29586), .A(n22726), .S(n21186), .Y(n29587) );
  MUX2X1 U19570 ( .B(n29592), .A(n29587), .S(n30281), .Y(n2249) );
  AOI22X1 U19571 ( .A(n29629), .B(n27321), .C(n29595), .D(n27317), .Y(n29589)
         );
  AOI22X1 U19572 ( .A(n34503), .B(n34197), .C(n29628), .D(n27320), .Y(n29588)
         );
  MUX2X1 U19573 ( .B(n25005), .A(n27181), .S(n30281), .Y(n29591) );
  AOI21X1 U19574 ( .A(loc_s2[5]), .B(n33993), .C(n24982), .Y(n29593) );
  AOI22X1 U19575 ( .A(n26339), .B(n24329), .C(n26274), .D(n29595), .Y(n29599)
         );
  AOI22X1 U19576 ( .A(n25721), .B(n29628), .C(n25715), .D(n34503), .Y(n29597)
         );
  NAND3X1 U19577 ( .A(n22282), .B(n24444), .C(n22734), .Y(n2250) );
  NAND3X1 U19578 ( .A(n25100), .B(wS), .C(n22939), .Y(n29623) );
  NAND3X1 U19579 ( .A(n20955), .B(net149749), .C(n29601), .Y(net90052) );
  AOI22X1 U19580 ( .A(n32191), .B(n27304), .C(n23443), .D(n15194), .Y(n29621)
         );
  NOR3X1 U19581 ( .A(oc[12]), .B(oc[16]), .C(n25702), .Y(n29611) );
  NOR3X1 U19582 ( .A(oc[30]), .B(oc[10]), .C(oc[8]), .Y(n29610) );
  NAND3X1 U19583 ( .A(n29611), .B(n29610), .C(n26069), .Y(n29727) );
  NOR3X1 U19584 ( .A(oc[11]), .B(oc[15]), .C(oc[13]), .Y(n29619) );
  NOR3X1 U19585 ( .A(oc[29]), .B(oc[9]), .C(oc[7]), .Y(n29618) );
  NOR3X1 U19586 ( .A(n24878), .B(addrLock), .C(net145105), .Y(n29622) );
  AOI21X1 U19587 ( .A(n23280), .B(n24246), .C(n29622), .Y(n29635) );
  NOR3X1 U19588 ( .A(n13801), .B(n13800), .C(n22979), .Y(n29625) );
  NAND3X1 U19589 ( .A(n29627), .B(n29626), .C(n29625), .Y(n30485) );
  AOI22X1 U19590 ( .A(n29629), .B(n25323), .C(n29628), .D(n25722), .Y(n29632)
         );
  AOI21X1 U19591 ( .A(n25715), .B(n29207), .C(n27300), .Y(n29630) );
  OAI21X1 U19592 ( .A(n34503), .B(n25447), .C(n23785), .Y(n29631) );
  OAI21X1 U19593 ( .A(Setup[1]), .B(n29703), .C(n27153), .Y(n33933) );
  AOI22X1 U19594 ( .A(n21055), .B(net114546), .C(net137830), .D(n33933), .Y(
        n29634) );
  OAI21X1 U19595 ( .A(n34385), .B(n23441), .C(n27113), .Y(n16195) );
  AOI21X1 U19596 ( .A(n29638), .B(n16187), .C(n16196), .Y(n29636) );
  OAI21X1 U19597 ( .A(n16195), .B(n26668), .C(n27113), .Y(n16242) );
  OAI21X1 U19598 ( .A(n27197), .B(n16196), .C(n27101), .Y(n29649) );
  XOR2X1 U19599 ( .A(n34501), .B(n34502), .Y(n16247) );
  OAI21X1 U19600 ( .A(n27100), .B(n16198), .C(n27193), .Y(n29637) );
  NOR3X1 U19601 ( .A(n29637), .B(n16242), .C(n34502), .Y(n34587) );
  XOR2X1 U19602 ( .A(n26803), .B(n34590), .Y(n16245) );
  XOR2X1 U19603 ( .A(n16187), .B(n29638), .Y(n16243) );
  XOR2X1 U19604 ( .A(n26812), .B(n29656), .Y(n16236) );
  XOR2X1 U19605 ( .A(n26339), .B(T[5]), .Y(n29648) );
  OAI21X1 U19606 ( .A(n26938), .B(n26812), .C(n26871), .Y(n29639) );
  OAI21X1 U19607 ( .A(T[5]), .B(n30186), .C(n26664), .Y(n16233) );
  XOR2X1 U19608 ( .A(n29655), .B(n29642), .Y(n16234) );
  OAI21X1 U19609 ( .A(n26938), .B(n29644), .C(n26871), .Y(n29646) );
  OAI21X1 U19610 ( .A(n26805), .B(n29643), .C(n26753), .Y(n29645) );
  MUX2X1 U19611 ( .B(n29646), .A(n29645), .S(n16233), .Y(n29647) );
  XOR2X1 U19612 ( .A(n26998), .B(n30281), .Y(n29651) );
  OAI21X1 U19613 ( .A(n26866), .B(n16213), .C(n26929), .Y(n16224) );
  OAI21X1 U19614 ( .A(n30186), .B(n29652), .C(n27162), .Y(n29653) );
  OAI21X1 U19615 ( .A(n34351), .B(n29653), .C(n26852), .Y(n16211) );
  NAND3X1 U19616 ( .A(n30410), .B(n21183), .C(n25447), .Y(n29657) );
  XOR2X1 U19617 ( .A(n24924), .B(n30281), .Y(n29659) );
  OAI21X1 U19618 ( .A(n25208), .B(n16132), .C(n26867), .Y(n16143) );
  OAI21X1 U19619 ( .A(n34351), .B(n27171), .C(n24965), .Y(n16130) );
  XOR2X1 U19620 ( .A(n25168), .B(n29683), .Y(n29666) );
  OAI21X1 U19621 ( .A(n29683), .B(n25168), .C(n23441), .Y(n29663) );
  OAI21X1 U19622 ( .A(n34385), .B(n25109), .C(n25207), .Y(n16114) );
  OAI21X1 U19623 ( .A(n25341), .B(n16115), .C(n25113), .Y(n29668) );
  XOR2X1 U19624 ( .A(n24938), .B(n30281), .Y(n29671) );
  OAI21X1 U19625 ( .A(n26928), .B(n16055), .C(n27076), .Y(n16066) );
  OAI21X1 U19626 ( .A(n34351), .B(n27075), .C(n24966), .Y(n16053) );
  NAND3X1 U19627 ( .A(n26163), .B(n20977), .C(n31917), .Y(n29678) );
  XOR2X1 U19628 ( .A(n25153), .B(n30281), .Y(n29677) );
  OAI21X1 U19629 ( .A(n25209), .B(n15981), .C(n26995), .Y(n15992) );
  OAI21X1 U19630 ( .A(n30186), .B(n25152), .C(n27162), .Y(n29681) );
  OAI21X1 U19631 ( .A(n34351), .B(n29681), .C(n26914), .Y(n15979) );
  XOR2X1 U19632 ( .A(n27098), .B(n29683), .Y(n29688) );
  AOI21X1 U19633 ( .A(n27098), .B(n23441), .C(n27301), .Y(n29684) );
  OAI21X1 U19634 ( .A(n25715), .B(n27176), .C(n23786), .Y(n29686) );
  OAI21X1 U19635 ( .A(n34385), .B(n29686), .C(n26994), .Y(n15963) );
  OAI21X1 U19636 ( .A(n26999), .B(n15964), .C(n26851), .Y(n29690) );
  NAND3X1 U19637 ( .A(n25489), .B(n34170), .C(n24867), .Y(n29694) );
  MUX2X1 U19638 ( .B(n24283), .A(n24323), .S(direct[0]), .Y(n29692) );
  MUX2X1 U19639 ( .B(n29692), .A(n15915), .S(direct[1]), .Y(n29693) );
  NAND3X1 U19640 ( .A(n24171), .B(n25778), .C(n29693), .Y(n29695) );
  OAI21X1 U19641 ( .A(n34172), .B(n29696), .C(net114546), .Y(n29702) );
  NAND3X1 U19642 ( .A(net110320), .B(net150385), .C(n27065), .Y(n29699) );
  NAND3X1 U19643 ( .A(n20818), .B(n24441), .C(net104600), .Y(n29700) );
  OAI21X1 U19644 ( .A(n34498), .B(n34555), .C(net64168), .Y(n29701) );
  NAND3X1 U19645 ( .A(n25072), .B(n29702), .C(n29701), .Y(n15900) );
  NAND3X1 U19646 ( .A(start), .B(net137830), .C(n29703), .Y(n29705) );
  NAND3X1 U19647 ( .A(oc[1]), .B(n29745), .C(n29755), .Y(n30001) );
  NAND3X1 U19648 ( .A(oc[23]), .B(oc[25]), .C(oc[27]), .Y(n29708) );
  NAND3X1 U19649 ( .A(oc[17]), .B(oc[21]), .C(oc[19]), .Y(n29707) );
  NOR3X1 U19650 ( .A(n24879), .B(n24889), .C(n23204), .Y(n29712) );
  NAND3X1 U19651 ( .A(oc[11]), .B(oc[15]), .C(oc[13]), .Y(n29710) );
  NAND3X1 U19652 ( .A(oc[29]), .B(oc[9]), .C(oc[7]), .Y(n29709) );
  AND2X2 U19653 ( .A(n29712), .B(n23745), .Y(n29947) );
  NAND3X1 U19654 ( .A(oc[5]), .B(n29713), .C(n29947), .Y(n29714) );
  NAND3X1 U19655 ( .A(oc[6]), .B(n21116), .C(n29715), .Y(n29721) );
  NAND3X1 U19656 ( .A(oc[24]), .B(oc[28]), .C(oc[26]), .Y(n29717) );
  NAND3X1 U19657 ( .A(oc[22]), .B(oc[20]), .C(oc[18]), .Y(n29716) );
  NAND3X1 U19658 ( .A(n25579), .B(n29946), .C(n23114), .Y(n29722) );
  NAND3X1 U19659 ( .A(n21224), .B(n25692), .C(n29756), .Y(n30036) );
  NOR3X1 U19660 ( .A(n29725), .B(n27059), .C(n23204), .Y(n29728) );
  OAI21X1 U19661 ( .A(n29978), .B(n27202), .C(n29215), .Y(n29729) );
  OAI21X1 U19662 ( .A(n21055), .B(n29732), .C(n29738), .Y(n29731) );
  AOI22X1 U19663 ( .A(n29352), .B(n29731), .C(n29750), .D(n27252), .Y(n29734)
         );
  OAI21X1 U19664 ( .A(n30556), .B(n25081), .C(n27208), .Y(n29733) );
  AOI21X1 U19665 ( .A(n27252), .B(n29331), .C(n33908), .Y(n29736) );
  OAI21X1 U19666 ( .A(n26735), .B(n27114), .C(n27273), .Y(n15873) );
  NAND3X1 U19667 ( .A(n30021), .B(n27252), .C(n29748), .Y(n29737) );
  OAI21X1 U19668 ( .A(n29738), .B(n29353), .C(n23787), .Y(n29743) );
  AOI21X1 U19669 ( .A(n30021), .B(n33908), .C(n29743), .Y(n29739) );
  OAI21X1 U19670 ( .A(n30062), .B(n25356), .C(n23788), .Y(n15880) );
  NAND3X1 U19671 ( .A(n21224), .B(oc[1]), .C(n29755), .Y(n29956) );
  NAND3X1 U19672 ( .A(n25107), .B(n24445), .C(n29740), .Y(n29742) );
  OAI21X1 U19673 ( .A(n29743), .B(n24685), .C(n14097), .Y(n15872) );
  NAND3X1 U19674 ( .A(oc[0]), .B(n29745), .C(n29756), .Y(n29989) );
  AOI22X1 U19675 ( .A(n29744), .B(n23285), .C(n22942), .D(n30038), .Y(n29747)
         );
  AOI21X1 U19676 ( .A(n29891), .B(n23285), .C(n29213), .Y(n29749) );
  OAI21X1 U19677 ( .A(n26880), .B(n27202), .C(n23789), .Y(n30489) );
  AOI21X1 U19678 ( .A(n27273), .B(n24993), .C(n29751), .Y(n29752) );
  NOR3X1 U19679 ( .A(n24888), .B(n29754), .C(n24892), .Y(n15865) );
  OAI21X1 U19680 ( .A(n30062), .B(n26820), .C(n26747), .Y(n29759) );
  NAND3X1 U19681 ( .A(n21224), .B(n21136), .C(n29755), .Y(n30023) );
  OAI21X1 U19682 ( .A(n33884), .B(n27217), .C(n30038), .Y(n29757) );
  OAI21X1 U19683 ( .A(n25332), .B(n26837), .C(n30491), .Y(n29758) );
  OAI21X1 U19684 ( .A(n29759), .B(n29758), .C(n14097), .Y(n15856) );
  AOI22X1 U19685 ( .A(n29744), .B(n23288), .C(n24928), .D(n30038), .Y(n29761)
         );
  OAI21X1 U19686 ( .A(n23287), .B(n26837), .C(n23749), .Y(n29764) );
  AOI21X1 U19687 ( .A(n29891), .B(n23288), .C(n29213), .Y(n29762) );
  OAI21X1 U19688 ( .A(n27016), .B(n27202), .C(n23790), .Y(n30494) );
  AOI21X1 U19689 ( .A(n27273), .B(n24995), .C(n29751), .Y(n29763) );
  NOR3X1 U19690 ( .A(n29764), .B(n29765), .C(n24893), .Y(n15844) );
  OAI21X1 U19691 ( .A(n30062), .B(n27103), .C(n26907), .Y(n29769) );
  OAI21X1 U19692 ( .A(n27205), .B(n26837), .C(n30496), .Y(n29768) );
  OAI21X1 U19693 ( .A(n29769), .B(n29768), .C(n14097), .Y(n15835) );
  AOI22X1 U19694 ( .A(n29744), .B(n23290), .C(n30038), .D(n27079), .Y(n29770)
         );
  OAI21X1 U19695 ( .A(n30495), .B(n26837), .C(n23750), .Y(n29773) );
  AOI21X1 U19696 ( .A(n29891), .B(n23290), .C(n29213), .Y(n29771) );
  OAI21X1 U19697 ( .A(n26821), .B(n27202), .C(n23791), .Y(n30499) );
  AOI21X1 U19698 ( .A(n27273), .B(n25123), .C(n29751), .Y(n29772) );
  NOR3X1 U19699 ( .A(n29773), .B(n29774), .C(n24894), .Y(n15823) );
  OAI21X1 U19700 ( .A(n30062), .B(n21375), .C(n24967), .Y(n29777) );
  OAI21X1 U19701 ( .A(n25830), .B(n27216), .C(n30038), .Y(n29775) );
  OAI21X1 U19702 ( .A(n32773), .B(n26837), .C(n30500), .Y(n29776) );
  OAI21X1 U19703 ( .A(n29777), .B(n29776), .C(n14097), .Y(n15814) );
  AOI22X1 U19704 ( .A(n29744), .B(n23293), .C(n23614), .D(n30038), .Y(n29778)
         );
  OAI21X1 U19705 ( .A(n23292), .B(n26837), .C(n23751), .Y(n29781) );
  AOI21X1 U19706 ( .A(n29891), .B(n23293), .C(n29213), .Y(n29779) );
  OAI21X1 U19707 ( .A(n26822), .B(n27202), .C(n23792), .Y(n30503) );
  AOI21X1 U19708 ( .A(n27273), .B(n24998), .C(n29751), .Y(n29780) );
  NOR3X1 U19709 ( .A(n29781), .B(n29782), .C(n24895), .Y(n15802) );
  OAI21X1 U19710 ( .A(n30062), .B(n27021), .C(n24968), .Y(n29785) );
  OAI21X1 U19711 ( .A(n33815), .B(n27219), .C(n30038), .Y(n29783) );
  OAI21X1 U19712 ( .A(n27119), .B(n26837), .C(n30505), .Y(n29784) );
  OAI21X1 U19713 ( .A(n29785), .B(n29784), .C(n14097), .Y(n15793) );
  AOI22X1 U19714 ( .A(n29744), .B(n23295), .C(n30038), .D(n26997), .Y(n29786)
         );
  OAI21X1 U19715 ( .A(n30504), .B(n26837), .C(n23752), .Y(n29789) );
  AOI21X1 U19716 ( .A(n29891), .B(n23295), .C(n29213), .Y(n29787) );
  OAI21X1 U19717 ( .A(n27017), .B(n27202), .C(n23793), .Y(n30508) );
  AOI21X1 U19718 ( .A(n27273), .B(n24999), .C(n29751), .Y(n29788) );
  NOR3X1 U19719 ( .A(n29789), .B(n29790), .C(n24896), .Y(n15781) );
  OAI21X1 U19720 ( .A(n30062), .B(n27191), .C(n26618), .Y(n29793) );
  OAI21X1 U19721 ( .A(n25771), .B(n27220), .C(n30038), .Y(n29791) );
  OAI21X1 U19722 ( .A(n27080), .B(n26837), .C(n30510), .Y(n29792) );
  OAI21X1 U19723 ( .A(n29793), .B(n29792), .C(n14097), .Y(n15772) );
  AOI22X1 U19724 ( .A(n29744), .B(n23298), .C(n30038), .D(n27174), .Y(n29795)
         );
  OAI21X1 U19725 ( .A(n30509), .B(n26837), .C(n23753), .Y(n29798) );
  AOI21X1 U19726 ( .A(n29891), .B(n23298), .C(n29213), .Y(n29796) );
  OAI21X1 U19727 ( .A(n26939), .B(n27202), .C(n23794), .Y(n30513) );
  AOI21X1 U19728 ( .A(n27273), .B(n25000), .C(n29751), .Y(n29797) );
  NOR3X1 U19729 ( .A(n29798), .B(n29799), .C(n24897), .Y(n15760) );
  OAI21X1 U19730 ( .A(n30062), .B(n21378), .C(n26644), .Y(n29802) );
  OAI21X1 U19731 ( .A(n23466), .B(n32988), .C(n30038), .Y(n29800) );
  OAI21X1 U19732 ( .A(n25770), .B(n26837), .C(n30515), .Y(n29801) );
  OAI21X1 U19733 ( .A(n29802), .B(n29801), .C(n14097), .Y(n15751) );
  AOI22X1 U19734 ( .A(n29744), .B(n29807), .C(n22943), .D(n30038), .Y(n29804)
         );
  OAI21X1 U19735 ( .A(n30514), .B(n26837), .C(n23754), .Y(n29809) );
  AOI21X1 U19736 ( .A(n29891), .B(n29807), .C(n29213), .Y(n29805) );
  OAI21X1 U19737 ( .A(n27082), .B(n27202), .C(n23795), .Y(n30518) );
  AOI21X1 U19738 ( .A(n27273), .B(n27061), .C(n29751), .Y(n29808) );
  NOR3X1 U19739 ( .A(n29809), .B(n29810), .C(n24898), .Y(n15738) );
  OAI21X1 U19740 ( .A(n30062), .B(n23111), .C(n24969), .Y(n29814) );
  OAI21X1 U19741 ( .A(n33748), .B(n21139), .C(n30038), .Y(n29812) );
  OAI21X1 U19742 ( .A(n27025), .B(n26837), .C(n30520), .Y(n29813) );
  OAI21X1 U19743 ( .A(n29814), .B(n29813), .C(n14097), .Y(n15729) );
  AOI22X1 U19744 ( .A(n29744), .B(n23299), .C(n22944), .D(n30038), .Y(n29816)
         );
  OAI21X1 U19745 ( .A(n30519), .B(n26837), .C(n23755), .Y(n29819) );
  AOI21X1 U19746 ( .A(n29891), .B(n23299), .C(n29213), .Y(n29817) );
  OAI21X1 U19747 ( .A(n29978), .B(n27116), .C(n23796), .Y(n30523) );
  AOI21X1 U19748 ( .A(n27273), .B(n25001), .C(n29751), .Y(n29818) );
  NOR3X1 U19749 ( .A(n29819), .B(n29820), .C(n24899), .Y(n15716) );
  OAI21X1 U19750 ( .A(n30062), .B(n26765), .C(n24970), .Y(n29823) );
  OAI21X1 U19751 ( .A(n26060), .B(n21188), .C(n30038), .Y(n29821) );
  OAI21X1 U19752 ( .A(n25147), .B(n26837), .C(n30524), .Y(n29822) );
  OAI21X1 U19753 ( .A(n29823), .B(n29822), .C(n14097), .Y(n15707) );
  AOI22X1 U19754 ( .A(n29744), .B(n23301), .C(n24929), .D(n30038), .Y(n29826)
         );
  OAI21X1 U19755 ( .A(n23300), .B(n26837), .C(n23756), .Y(n29829) );
  AOI21X1 U19756 ( .A(n29891), .B(n23301), .C(n29213), .Y(n29827) );
  OAI21X1 U19757 ( .A(n26880), .B(n27116), .C(n23797), .Y(n30527) );
  AOI21X1 U19758 ( .A(n27273), .B(n25161), .C(n29751), .Y(n29828) );
  NOR3X1 U19759 ( .A(n29829), .B(n29830), .C(n24900), .Y(n15695) );
  OAI21X1 U19760 ( .A(n30062), .B(n26942), .C(n24971), .Y(n29834) );
  OAI21X1 U19761 ( .A(n23468), .B(n21178), .C(n30038), .Y(n29832) );
  OAI21X1 U19762 ( .A(n25148), .B(n26837), .C(n30528), .Y(n29833) );
  OAI21X1 U19763 ( .A(n29834), .B(n29833), .C(n14097), .Y(n15686) );
  AOI22X1 U19764 ( .A(n29744), .B(n23282), .C(n24930), .D(n30038), .Y(n29837)
         );
  OAI21X1 U19765 ( .A(n23302), .B(n26837), .C(n23757), .Y(n29840) );
  AOI21X1 U19766 ( .A(n29891), .B(n23282), .C(n29213), .Y(n29838) );
  OAI21X1 U19767 ( .A(n27016), .B(n27116), .C(n23798), .Y(n30531) );
  AOI21X1 U19768 ( .A(n27273), .B(n24992), .C(n29751), .Y(n29839) );
  NOR3X1 U19769 ( .A(n29840), .B(n29841), .C(n24901), .Y(n15674) );
  OAI21X1 U19770 ( .A(n30062), .B(n33682), .C(n26676), .Y(n29844) );
  OAI21X1 U19771 ( .A(n23469), .B(n27232), .C(n30038), .Y(n29842) );
  OAI21X1 U19772 ( .A(n25149), .B(n26837), .C(n30532), .Y(n29843) );
  OAI21X1 U19773 ( .A(n29844), .B(n29843), .C(n14097), .Y(n15665) );
  NAND3X1 U19774 ( .A(n29845), .B(oc[5]), .C(n23113), .Y(n32971) );
  AOI22X1 U19775 ( .A(n29744), .B(n23283), .C(n24931), .D(n30038), .Y(n29847)
         );
  OAI21X1 U19776 ( .A(n23303), .B(n26837), .C(n23758), .Y(n29850) );
  AOI21X1 U19777 ( .A(n29891), .B(n23283), .C(n29213), .Y(n29848) );
  OAI21X1 U19778 ( .A(n26821), .B(n27116), .C(n23799), .Y(n30535) );
  AOI21X1 U19779 ( .A(n27273), .B(n25120), .C(n29751), .Y(n29849) );
  NOR3X1 U19780 ( .A(n29850), .B(n29851), .C(n24902), .Y(n15653) );
  OAI21X1 U19781 ( .A(n30062), .B(n27207), .C(n26707), .Y(n29854) );
  OAI21X1 U19782 ( .A(n26519), .B(n21220), .C(n30038), .Y(n29852) );
  OAI21X1 U19783 ( .A(n32953), .B(n26837), .C(n30537), .Y(n29853) );
  OAI21X1 U19784 ( .A(n29854), .B(n29853), .C(n14097), .Y(n15644) );
  AOI22X1 U19785 ( .A(n29744), .B(n23286), .C(n22945), .D(n30038), .Y(n29855)
         );
  OAI21X1 U19786 ( .A(n30536), .B(n26837), .C(n23759), .Y(n29858) );
  AOI21X1 U19787 ( .A(n29891), .B(n23286), .C(n29213), .Y(n29856) );
  OAI21X1 U19788 ( .A(n26822), .B(n27116), .C(n23800), .Y(n30540) );
  AOI21X1 U19789 ( .A(n27273), .B(n24994), .C(n29751), .Y(n29857) );
  NOR3X1 U19790 ( .A(n29858), .B(n29859), .C(n24903), .Y(n15632) );
  OAI21X1 U19791 ( .A(n30062), .B(n25440), .C(n24972), .Y(n29862) );
  OAI21X1 U19792 ( .A(n33639), .B(n21152), .C(n30038), .Y(n29860) );
  OAI21X1 U19793 ( .A(n27023), .B(n26837), .C(n30542), .Y(n29861) );
  OAI21X1 U19794 ( .A(n29862), .B(n29861), .C(n14097), .Y(n15623) );
  AOI22X1 U19795 ( .A(n29744), .B(n23289), .C(n22946), .D(n30038), .Y(n29863)
         );
  OAI21X1 U19796 ( .A(n30541), .B(n26837), .C(n23760), .Y(n29866) );
  AOI21X1 U19797 ( .A(n29891), .B(n23289), .C(n29213), .Y(n29864) );
  OAI21X1 U19798 ( .A(n27017), .B(n27116), .C(n23801), .Y(n30545) );
  AOI21X1 U19799 ( .A(n27273), .B(n24996), .C(n29751), .Y(n29865) );
  NOR3X1 U19800 ( .A(n29866), .B(n29867), .C(n24904), .Y(n15611) );
  OAI21X1 U19801 ( .A(n30062), .B(n26940), .C(n26748), .Y(n29870) );
  OAI21X1 U19802 ( .A(n26518), .B(n27225), .C(n30038), .Y(n29868) );
  OAI21X1 U19803 ( .A(n22948), .B(n26837), .C(n30547), .Y(n29869) );
  OAI21X1 U19804 ( .A(n29870), .B(n29869), .C(n14097), .Y(n15601) );
  AOI22X1 U19805 ( .A(n29744), .B(n23291), .C(n22949), .D(n30038), .Y(n29872)
         );
  OAI21X1 U19806 ( .A(n30546), .B(n26837), .C(n23761), .Y(n29875) );
  AOI21X1 U19807 ( .A(n29891), .B(n23291), .C(n29213), .Y(n29873) );
  OAI21X1 U19808 ( .A(n26939), .B(n27116), .C(n23802), .Y(n30550) );
  AOI21X1 U19809 ( .A(n27273), .B(n24997), .C(n29751), .Y(n29874) );
  NOR3X1 U19810 ( .A(n29875), .B(n27275), .C(n24905), .Y(n15589) );
  AOI21X1 U19811 ( .A(n30038), .B(n24248), .C(n30556), .Y(n30551) );
  AOI21X1 U19812 ( .A(n30038), .B(n33587), .C(n27275), .Y(n29877) );
  NAND3X1 U19813 ( .A(n25106), .B(n25117), .C(n24847), .Y(n29878) );
  NAND2X1 U19814 ( .A(n14097), .B(n23905), .Y(n15574) );
  NAND3X1 U19815 ( .A(n33558), .B(n27273), .C(n26078), .Y(n29884) );
  AOI21X1 U19816 ( .A(n29879), .B(n29967), .C(n29213), .Y(n29880) );
  OAI21X1 U19817 ( .A(n25002), .B(n26932), .C(n23803), .Y(n33555) );
  OAI21X1 U19818 ( .A(n29882), .B(n29353), .C(n25117), .Y(n29883) );
  AOI21X1 U19819 ( .A(n24257), .B(n27208), .C(n29883), .Y(n15566) );
  OAI21X1 U19820 ( .A(n29886), .B(n27114), .C(n27273), .Y(n29885) );
  OAI21X1 U19821 ( .A(n27249), .B(n33555), .C(n29352), .Y(n29888) );
  AOI22X1 U19822 ( .A(n29750), .B(n23294), .C(n29744), .D(n23294), .Y(n29887)
         );
  NAND3X1 U19823 ( .A(n29894), .B(n29888), .C(n24697), .Y(n29889) );
  AOI21X1 U19824 ( .A(n29966), .B(n21211), .C(n29213), .Y(n29890) );
  OAI21X1 U19825 ( .A(n25128), .B(n26932), .C(n23804), .Y(n30557) );
  OAI21X1 U19826 ( .A(n27249), .B(n30557), .C(n29352), .Y(n29893) );
  AOI22X1 U19827 ( .A(n29750), .B(n23296), .C(n29744), .D(n23296), .Y(n29892)
         );
  NAND3X1 U19828 ( .A(n29894), .B(n29893), .C(n24698), .Y(n29895) );
  NAND3X1 U19829 ( .A(n30555), .B(n27273), .C(n25403), .Y(n29899) );
  OAI21X1 U19830 ( .A(n29897), .B(n29353), .C(n23889), .Y(n29898) );
  AOI21X1 U19831 ( .A(n24258), .B(n27208), .C(n29898), .Y(n15535) );
  AOI22X1 U19832 ( .A(n29744), .B(n29902), .C(n22951), .D(n30038), .Y(n29900)
         );
  OAI21X1 U19833 ( .A(n30558), .B(n26837), .C(n23762), .Y(n29904) );
  AOI21X1 U19834 ( .A(n29891), .B(n29902), .C(n29213), .Y(n29901) );
  OAI21X1 U19835 ( .A(n26880), .B(n27201), .C(n23805), .Y(n30562) );
  AOI21X1 U19836 ( .A(n27273), .B(n26853), .C(n29751), .Y(n29903) );
  NOR3X1 U19837 ( .A(n29904), .B(n29907), .C(n24906), .Y(n15521) );
  OAI21X1 U19838 ( .A(n33531), .B(n30556), .C(n27208), .Y(n29908) );
  AOI22X1 U19839 ( .A(n30021), .B(n24303), .C(n30038), .D(n25134), .Y(n29906)
         );
  NAND3X1 U19840 ( .A(n29908), .B(n26794), .C(n24699), .Y(n29909) );
  NAND2X1 U19841 ( .A(n14097), .B(n23906), .Y(n15512) );
  AOI22X1 U19842 ( .A(n29744), .B(n30033), .C(n23633), .D(n30038), .Y(n29910)
         );
  OAI21X1 U19843 ( .A(n23273), .B(n26837), .C(n23763), .Y(n29914) );
  AOI21X1 U19844 ( .A(n29891), .B(n30033), .C(n29213), .Y(n29911) );
  OAI21X1 U19845 ( .A(n27016), .B(n27201), .C(n23806), .Y(n30566) );
  AOI21X1 U19846 ( .A(n27273), .B(n26798), .C(n29751), .Y(n29913) );
  NOR3X1 U19847 ( .A(n29914), .B(n29917), .C(n24907), .Y(n15500) );
  OAI21X1 U19848 ( .A(n33508), .B(n30556), .C(n27208), .Y(n29918) );
  AOI22X1 U19849 ( .A(n30021), .B(n24304), .C(n30038), .D(n25135), .Y(n29916)
         );
  NAND3X1 U19850 ( .A(n29918), .B(n26912), .C(n24700), .Y(n29919) );
  NAND2X1 U19851 ( .A(n14097), .B(n23907), .Y(n15490) );
  AOI22X1 U19852 ( .A(n29744), .B(n29922), .C(n22952), .D(n30038), .Y(n29920)
         );
  OAI21X1 U19853 ( .A(n30567), .B(n26837), .C(n23764), .Y(n29924) );
  AOI21X1 U19854 ( .A(n29891), .B(n29922), .C(n29213), .Y(n29921) );
  OAI21X1 U19855 ( .A(n26821), .B(n27201), .C(n23807), .Y(n30571) );
  AOI21X1 U19856 ( .A(n27273), .B(n26752), .C(n29751), .Y(n29923) );
  NOR3X1 U19857 ( .A(n29924), .B(n29928), .C(n24908), .Y(n15478) );
  OAI21X1 U19858 ( .A(n33485), .B(n30556), .C(n27208), .Y(n29929) );
  AOI22X1 U19859 ( .A(n30021), .B(n24305), .C(n30038), .D(n25136), .Y(n29927)
         );
  NAND3X1 U19860 ( .A(n29929), .B(n25073), .C(n24701), .Y(n29930) );
  NAND2X1 U19861 ( .A(n14097), .B(n23908), .Y(n15469) );
  AOI22X1 U19862 ( .A(n29744), .B(n29933), .C(n22953), .D(n30038), .Y(n29931)
         );
  OAI21X1 U19863 ( .A(n30572), .B(n26837), .C(n23765), .Y(n29935) );
  AOI21X1 U19864 ( .A(n29891), .B(n29933), .C(n29213), .Y(n29932) );
  OAI21X1 U19865 ( .A(n26822), .B(n27201), .C(n23808), .Y(n30576) );
  AOI21X1 U19866 ( .A(n27273), .B(n26710), .C(n29751), .Y(n29934) );
  NOR3X1 U19867 ( .A(n29935), .B(n29938), .C(n24909), .Y(n15456) );
  OAI21X1 U19868 ( .A(n33462), .B(n30556), .C(n27208), .Y(n29939) );
  NAND3X1 U19869 ( .A(n29967), .B(n27315), .C(n21106), .Y(n32529) );
  AOI22X1 U19870 ( .A(n30021), .B(n24306), .C(n30038), .D(n25137), .Y(n29937)
         );
  NAND3X1 U19871 ( .A(n29939), .B(n25074), .C(n24702), .Y(n29940) );
  NAND2X1 U19872 ( .A(n14097), .B(n23909), .Y(n15446) );
  AOI22X1 U19873 ( .A(n29744), .B(n29943), .C(n22954), .D(n30038), .Y(n29941)
         );
  OAI21X1 U19874 ( .A(n30577), .B(n26837), .C(n23766), .Y(n29945) );
  AOI21X1 U19875 ( .A(n29891), .B(n29943), .C(n29213), .Y(n29942) );
  OAI21X1 U19876 ( .A(n27017), .B(n27201), .C(n23809), .Y(n30581) );
  AOI21X1 U19877 ( .A(n27273), .B(n26983), .C(n29751), .Y(n29944) );
  NOR3X1 U19878 ( .A(n29945), .B(n29951), .C(n24910), .Y(n15434) );
  OAI21X1 U19879 ( .A(n25774), .B(n30556), .C(n27208), .Y(n29952) );
  NAND3X1 U19880 ( .A(oc[6]), .B(n29946), .C(n29947), .Y(n29948) );
  AOI22X1 U19881 ( .A(n30021), .B(n24307), .C(n30038), .D(n25138), .Y(n29950)
         );
  NAND3X1 U19882 ( .A(n29952), .B(n26848), .C(n24703), .Y(n29953) );
  NAND2X1 U19883 ( .A(n14097), .B(n23910), .Y(n15424) );
  AOI22X1 U19884 ( .A(n29744), .B(n23284), .C(n22955), .D(n30038), .Y(n29954)
         );
  OAI21X1 U19885 ( .A(n30582), .B(n26837), .C(n23767), .Y(n29958) );
  AOI21X1 U19886 ( .A(n29891), .B(n23444), .C(n29213), .Y(n29955) );
  OAI21X1 U19887 ( .A(n26939), .B(n27201), .C(n23810), .Y(n30586) );
  AOI21X1 U19888 ( .A(n27273), .B(n25121), .C(n29751), .Y(n29957) );
  NOR3X1 U19889 ( .A(n29958), .B(n29961), .C(n24911), .Y(n15411) );
  OAI21X1 U19890 ( .A(n33417), .B(n30556), .C(n27208), .Y(n29962) );
  AOI22X1 U19891 ( .A(n30021), .B(n24308), .C(n30038), .D(n25139), .Y(n29960)
         );
  NAND3X1 U19892 ( .A(n29962), .B(n26750), .C(n24704), .Y(n29963) );
  NAND2X1 U19893 ( .A(n14097), .B(n23911), .Y(n15401) );
  AOI22X1 U19894 ( .A(n29744), .B(n29968), .C(n22956), .D(n30038), .Y(n29964)
         );
  OAI21X1 U19895 ( .A(n30587), .B(n26837), .C(n23768), .Y(n29970) );
  AOI21X1 U19896 ( .A(n29891), .B(n29968), .C(n29213), .Y(n29965) );
  OAI21X1 U19897 ( .A(n27082), .B(n27201), .C(n23811), .Y(n30591) );
  AOI21X1 U19898 ( .A(n27273), .B(n26916), .C(n29751), .Y(n29969) );
  NOR3X1 U19899 ( .A(n29970), .B(n29973), .C(n24912), .Y(n15387) );
  OAI21X1 U19900 ( .A(n25657), .B(n30556), .C(n27208), .Y(n29974) );
  AOI22X1 U19901 ( .A(n30021), .B(n24309), .C(n30038), .D(n25140), .Y(n29972)
         );
  NAND3X1 U19902 ( .A(n29974), .B(n26979), .C(n24705), .Y(n29975) );
  NAND2X1 U19903 ( .A(n14097), .B(n23912), .Y(n15377) );
  AOI22X1 U19904 ( .A(n29744), .B(n23446), .C(n22957), .D(n30038), .Y(n29976)
         );
  OAI21X1 U19905 ( .A(n30592), .B(n26837), .C(n23769), .Y(n29981) );
  AOI21X1 U19906 ( .A(n29891), .B(n23446), .C(n29213), .Y(n29977) );
  OAI21X1 U19907 ( .A(n29978), .B(n26948), .C(n23812), .Y(n30596) );
  AOI21X1 U19908 ( .A(n27273), .B(n25122), .C(n29751), .Y(n29980) );
  NOR3X1 U19909 ( .A(n29981), .B(n29984), .C(n24913), .Y(n15362) );
  OAI21X1 U19910 ( .A(n25680), .B(n30556), .C(n27208), .Y(n29985) );
  AOI22X1 U19911 ( .A(n30021), .B(n24310), .C(n30038), .D(n25141), .Y(n29983)
         );
  NAND3X1 U19912 ( .A(n29985), .B(n25075), .C(n24706), .Y(n29986) );
  NAND2X1 U19913 ( .A(n14097), .B(n23913), .Y(n15352) );
  AOI22X1 U19914 ( .A(n29744), .B(n29993), .C(n22958), .D(n30038), .Y(n29987)
         );
  OAI21X1 U19915 ( .A(n30597), .B(n26837), .C(n23770), .Y(n29992) );
  AOI21X1 U19916 ( .A(n29891), .B(n29993), .C(n29213), .Y(n29988) );
  OAI21X1 U19917 ( .A(n26880), .B(n26948), .C(n23813), .Y(n30601) );
  AOI21X1 U19918 ( .A(n27273), .B(n25194), .C(n29751), .Y(n29991) );
  NOR3X1 U19919 ( .A(n29992), .B(n29996), .C(n24914), .Y(n15339) );
  OAI21X1 U19920 ( .A(n33326), .B(n30556), .C(n27208), .Y(n29997) );
  AOI22X1 U19921 ( .A(n30021), .B(n24311), .C(n30038), .D(n25142), .Y(n29995)
         );
  NAND3X1 U19922 ( .A(n29997), .B(n26795), .C(n24707), .Y(n29998) );
  NAND2X1 U19923 ( .A(n14097), .B(n23914), .Y(n15329) );
  AOI22X1 U19924 ( .A(n29744), .B(n30002), .C(n22959), .D(n30038), .Y(n29999)
         );
  OAI21X1 U19925 ( .A(n30602), .B(n26837), .C(n23771), .Y(n30004) );
  AOI21X1 U19926 ( .A(n29891), .B(n30002), .C(n29213), .Y(n30000) );
  OAI21X1 U19927 ( .A(n27016), .B(n26948), .C(n23814), .Y(n30606) );
  AOI21X1 U19928 ( .A(n27273), .B(n26984), .C(n29751), .Y(n30003) );
  NOR3X1 U19929 ( .A(n30004), .B(n30007), .C(n24915), .Y(n15316) );
  OAI21X1 U19930 ( .A(n33295), .B(n30556), .C(n27208), .Y(n30008) );
  AOI22X1 U19931 ( .A(n30021), .B(n24312), .C(n30038), .D(n25143), .Y(n30006)
         );
  NAND3X1 U19932 ( .A(n30008), .B(n26849), .C(n24708), .Y(n30009) );
  NAND2X1 U19933 ( .A(n14097), .B(n23915), .Y(n15306) );
  AOI22X1 U19934 ( .A(n29744), .B(n23447), .C(n22960), .D(n30038), .Y(n30010)
         );
  OAI21X1 U19935 ( .A(n30607), .B(n26837), .C(n23772), .Y(n30014) );
  AOI21X1 U19936 ( .A(n29891), .B(n23447), .C(n29214), .Y(n30011) );
  OAI21X1 U19937 ( .A(n26821), .B(n26948), .C(n23815), .Y(n30611) );
  AOI21X1 U19938 ( .A(n27273), .B(n25124), .C(n29751), .Y(n30013) );
  NOR3X1 U19939 ( .A(n30014), .B(n30017), .C(n24916), .Y(n15293) );
  OAI21X1 U19940 ( .A(n25658), .B(n30556), .C(n27208), .Y(n30018) );
  AOI22X1 U19941 ( .A(n30021), .B(n24313), .C(n30038), .D(n25144), .Y(n30016)
         );
  NAND3X1 U19942 ( .A(n30018), .B(n25076), .C(n24709), .Y(n30019) );
  NAND2X1 U19943 ( .A(n14097), .B(n23916), .Y(n15283) );
  AOI22X1 U19944 ( .A(n29744), .B(n23449), .C(n22961), .D(n30038), .Y(n30020)
         );
  OAI21X1 U19945 ( .A(n30612), .B(n26837), .C(n23773), .Y(n30026) );
  AOI21X1 U19946 ( .A(n29891), .B(n23448), .C(n29214), .Y(n30022) );
  OAI21X1 U19947 ( .A(n26822), .B(n26948), .C(n23816), .Y(n30618) );
  AOI21X1 U19948 ( .A(n27273), .B(n25125), .C(n29751), .Y(n30025) );
  NOR3X1 U19949 ( .A(n30026), .B(n30030), .C(n24917), .Y(n15269) );
  OAI21X1 U19950 ( .A(n33234), .B(n30556), .C(n27208), .Y(n30031) );
  AOI22X1 U19951 ( .A(n30021), .B(n24314), .C(n30038), .D(n25118), .Y(n30029)
         );
  NAND3X1 U19952 ( .A(n30031), .B(n25077), .C(n24710), .Y(n30032) );
  NAND2X1 U19953 ( .A(n14097), .B(n23917), .Y(n15260) );
  AOI21X1 U19954 ( .A(n29891), .B(n30040), .C(n29214), .Y(n30034) );
  OAI21X1 U19955 ( .A(n27017), .B(n26948), .C(n23817), .Y(n30037) );
  OAI21X1 U19956 ( .A(n21055), .B(n23308), .C(n30622), .Y(n30039) );
  OAI21X1 U19957 ( .A(n26879), .B(n27114), .C(n27273), .Y(n30617) );
  AOI21X1 U19958 ( .A(n29352), .B(n30039), .C(n30617), .Y(n30043) );
  OAI21X1 U19959 ( .A(n24279), .B(n26799), .C(n27195), .Y(n30041) );
  AOI22X1 U19960 ( .A(n30038), .B(n30041), .C(n29750), .D(n30040), .Y(n30042)
         );
  NAND3X1 U19961 ( .A(n8037), .B(n30045), .C(n30044), .Y(n30049) );
  AOI21X1 U19962 ( .A(n8034), .B(n30047), .C(n30046), .Y(n30048) );
  OAI21X1 U19963 ( .A(n25127), .B(n21093), .C(net125066), .Y(n30052) );
  AOI21X1 U19964 ( .A(net109585), .B(n30052), .C(n30051), .Y(n15222) );
  AOI21X1 U19965 ( .A(n21030), .B(n25663), .C(n24033), .Y(n30059) );
  AOI22X1 U19966 ( .A(n21117), .B(n25763), .C(locTrig[2]), .D(n25760), .Y(
        n30058) );
  OAI21X1 U19967 ( .A(net110411), .B(n30054), .C(n20818), .Y(n30055) );
  AOI21X1 U19968 ( .A(n21117), .B(n26062), .C(n30055), .Y(n30057) );
  AOI22X1 U19969 ( .A(locTrig[2]), .B(net109176), .C(locTrig[3]), .D(net108619), .Y(n30056) );
  AOI22X1 U19970 ( .A(n24325), .B(n24302), .C(n24694), .D(n24696), .Y(n30060)
         );
  OAI21X1 U19971 ( .A(n24271), .B(net108653), .C(n21432), .Y(n30063) );
  NOR3X1 U19972 ( .A(n30063), .B(n25211), .C(n25116), .Y(n15205) );
  NAND2X1 U19973 ( .A(n14097), .B(n23280), .Y(n15204) );
  NAND3X1 U19974 ( .A(n23443), .B(n30066), .C(n24869), .Y(n30069) );
  NAND3X1 U19975 ( .A(n24172), .B(n26056), .C(n24870), .Y(n15196) );
  OAI21X1 U19976 ( .A(n15183), .B(net110411), .C(n30070), .Y(n15189) );
  OAI21X1 U19977 ( .A(n15183), .B(n25836), .C(n30070), .Y(n15187) );
  OAI21X1 U19978 ( .A(n15183), .B(net94647), .C(n30070), .Y(n15185) );
  OAI21X1 U19979 ( .A(n15183), .B(net94645), .C(n30070), .Y(n15181) );
  NAND3X1 U19980 ( .A(n30327), .B(n30371), .C(n30234), .Y(n30071) );
  NAND3X1 U19981 ( .A(n30126), .B(n30117), .C(n30100), .Y(n30072) );
  AOI22X1 U19982 ( .A(n31916), .B(n29320), .C(n29441), .D(n25715), .Y(n30084)
         );
  OAI21X1 U19983 ( .A(Setup[1]), .B(net111600), .C(n24964), .Y(n30074) );
  NAND3X1 U19984 ( .A(n30643), .B(n29353), .C(n24871), .Y(n30471) );
  NAND3X1 U19985 ( .A(n30079), .B(n23443), .C(n21196), .Y(n30630) );
  AOI21X1 U19986 ( .A(n23311), .B(n34498), .C(n30080), .Y(n30081) );
  OAI21X1 U19987 ( .A(n25357), .B(n29219), .C(n23818), .Y(n30082) );
  AOI22X1 U19988 ( .A(n30080), .B(n29217), .C(net64168), .D(n30082), .Y(n30083) );
  NAND3X1 U19989 ( .A(data_in[0]), .B(n30117), .C(n30100), .Y(n30085) );
  AOI22X1 U19990 ( .A(n30670), .B(n29320), .C(n29440), .D(n32199), .Y(n30091)
         );
  AOI21X1 U19991 ( .A(n23312), .B(n34498), .C(n30087), .Y(n30088) );
  OAI21X1 U19992 ( .A(n26935), .B(n29219), .C(n23819), .Y(n30089) );
  AOI22X1 U19993 ( .A(n30087), .B(n29217), .C(net64168), .D(n30089), .Y(n30090) );
  NAND3X1 U19994 ( .A(data_in[1]), .B(n30126), .C(n30100), .Y(n30092) );
  AOI22X1 U19995 ( .A(n31927), .B(n29320), .C(n29441), .D(n32204), .Y(n30099)
         );
  NAND3X1 U19996 ( .A(n21089), .B(n21231), .C(n26505), .Y(n30093) );
  NAND3X1 U19997 ( .A(net149983), .B(net150133), .C(net105803), .Y(n30094) );
  AOI21X1 U19998 ( .A(n23313), .B(n34498), .C(n30095), .Y(n30096) );
  OAI21X1 U19999 ( .A(n27090), .B(n29219), .C(n23820), .Y(n30097) );
  AOI22X1 U20000 ( .A(n30095), .B(n29217), .C(net64168), .D(n30097), .Y(n30098) );
  NAND3X1 U20001 ( .A(data_in[0]), .B(data_in[1]), .C(n30100), .Y(n30101) );
  AOI22X1 U20002 ( .A(n30713), .B(n29320), .C(n29440), .D(n32209), .Y(n30108)
         );
  NAND3X1 U20003 ( .A(n26142), .B(n21231), .C(n26485), .Y(n30102) );
  NAND3X1 U20004 ( .A(net149983), .B(net150126), .C(net105808), .Y(n30103) );
  AOI21X1 U20005 ( .A(n23314), .B(n34498), .C(n30104), .Y(n30105) );
  OAI21X1 U20006 ( .A(n26816), .B(n29219), .C(n23821), .Y(n30106) );
  AOI22X1 U20007 ( .A(n30104), .B(n29217), .C(net64168), .D(n30106), .Y(n30107) );
  NAND3X1 U20008 ( .A(data_in[2]), .B(n30126), .C(n30117), .Y(n30109) );
  AOI22X1 U20009 ( .A(n31937), .B(n29320), .C(n29441), .D(n32214), .Y(n30116)
         );
  NAND3X1 U20010 ( .A(n21089), .B(n26514), .C(n28604), .Y(n30110) );
  NAND3X1 U20011 ( .A(net105821), .B(net150133), .C(net151834), .Y(n30111) );
  AOI21X1 U20012 ( .A(n23315), .B(n34498), .C(n30112), .Y(n30113) );
  OAI21X1 U20013 ( .A(n27088), .B(n29219), .C(n23822), .Y(n30114) );
  AOI22X1 U20014 ( .A(n30112), .B(n29217), .C(net64168), .D(n30114), .Y(n30115) );
  NAND3X1 U20015 ( .A(data_in[2]), .B(data_in[0]), .C(n30117), .Y(n30118) );
  AOI22X1 U20016 ( .A(n30753), .B(n29320), .C(n29440), .D(n32219), .Y(n30125)
         );
  NAND3X1 U20017 ( .A(n26143), .B(n26514), .C(n28605), .Y(n30119) );
  NAND3X1 U20018 ( .A(net105821), .B(net111222), .C(net149936), .Y(n30120) );
  AOI21X1 U20019 ( .A(n23316), .B(n34498), .C(n30121), .Y(n30122) );
  OAI21X1 U20020 ( .A(n26761), .B(n29219), .C(n23823), .Y(n30123) );
  AOI22X1 U20021 ( .A(n30121), .B(n29217), .C(net64168), .D(n30123), .Y(n30124) );
  AOI22X1 U20022 ( .A(n31947), .B(n29320), .C(n29441), .D(n32224), .Y(n30134)
         );
  NAND3X1 U20023 ( .A(n26517), .B(n28605), .C(n26485), .Y(n30128) );
  NAND3X1 U20024 ( .A(net149982), .B(net150133), .C(net105819), .Y(n30129) );
  AOI21X1 U20025 ( .A(n23317), .B(n34498), .C(n30130), .Y(n30131) );
  OAI21X1 U20026 ( .A(n27002), .B(n29219), .C(n23824), .Y(n30132) );
  AOI22X1 U20027 ( .A(n30130), .B(n29217), .C(net64168), .D(n30132), .Y(n30133) );
  AOI22X1 U20028 ( .A(n30793), .B(n29320), .C(n29440), .D(n32229), .Y(n30142)
         );
  NAND3X1 U20029 ( .A(n26087), .B(n28605), .C(n26507), .Y(n30136) );
  NAND3X1 U20030 ( .A(net113308), .B(net149936), .C(net105859), .Y(n30137) );
  INVX2 U20031 ( .A(n22675), .Y(n30473) );
  AOI21X1 U20032 ( .A(n31955), .B(n34498), .C(n30138), .Y(n30139) );
  OAI21X1 U20033 ( .A(n26875), .B(n29219), .C(n23825), .Y(n30140) );
  AOI22X1 U20034 ( .A(n30138), .B(n29217), .C(net64168), .D(n30140), .Y(n30141) );
  NAND3X1 U20035 ( .A(data_in[3]), .B(n30327), .C(n30234), .Y(n30143) );
  AOI22X1 U20036 ( .A(n31958), .B(n29320), .C(n29441), .D(n32234), .Y(n30148)
         );
  AOI21X1 U20037 ( .A(n23318), .B(n34498), .C(n30144), .Y(n30145) );
  OAI21X1 U20038 ( .A(n26716), .B(n29219), .C(n23826), .Y(n30146) );
  AOI22X1 U20039 ( .A(n30144), .B(n29217), .C(net64168), .D(n30146), .Y(n30147) );
  AOI22X1 U20040 ( .A(n30833), .B(n29320), .C(n29440), .D(n32239), .Y(n30153)
         );
  AOI21X1 U20041 ( .A(n23319), .B(n34498), .C(n30149), .Y(n30150) );
  OAI21X1 U20042 ( .A(n26763), .B(n29219), .C(n23827), .Y(n30151) );
  AOI22X1 U20043 ( .A(n30149), .B(n29217), .C(net64168), .D(n30151), .Y(n30152) );
  AOI22X1 U20044 ( .A(n31968), .B(n29320), .C(n29441), .D(n32244), .Y(n30158)
         );
  AOI21X1 U20045 ( .A(n23320), .B(n34498), .C(n30154), .Y(n30155) );
  OAI21X1 U20046 ( .A(n26937), .B(n29219), .C(n23828), .Y(n30156) );
  AOI22X1 U20047 ( .A(n30154), .B(n29217), .C(net64168), .D(n30156), .Y(n30157) );
  AOI22X1 U20048 ( .A(n30873), .B(n29320), .C(n29440), .D(n32249), .Y(n30163)
         );
  AOI21X1 U20049 ( .A(n23322), .B(n34498), .C(n30159), .Y(n30160) );
  OAI21X1 U20050 ( .A(n26877), .B(n29219), .C(n23829), .Y(n30161) );
  AOI22X1 U20051 ( .A(n30159), .B(n29217), .C(net64168), .D(n30161), .Y(n30162) );
  AOI22X1 U20052 ( .A(n31977), .B(n29320), .C(n29440), .D(n32254), .Y(n30168)
         );
  AOI21X1 U20053 ( .A(n23323), .B(n34498), .C(n30164), .Y(n30165) );
  OAI21X1 U20054 ( .A(n27004), .B(n29219), .C(n23830), .Y(n30166) );
  AOI22X1 U20055 ( .A(n30164), .B(n29217), .C(net64168), .D(n30166), .Y(n30167) );
  AOI22X1 U20056 ( .A(n30914), .B(n29320), .C(n29441), .D(n32259), .Y(n30173)
         );
  AOI21X1 U20057 ( .A(n23324), .B(n34498), .C(n30169), .Y(n30170) );
  OAI21X1 U20058 ( .A(n26818), .B(n29219), .C(n23831), .Y(n30171) );
  AOI22X1 U20059 ( .A(n30169), .B(n29217), .C(net64168), .D(n30171), .Y(n30172) );
  AOI22X1 U20060 ( .A(n31987), .B(n29320), .C(n29440), .D(n32264), .Y(n30178)
         );
  AOI21X1 U20061 ( .A(n32266), .B(n34498), .C(n30174), .Y(n30175) );
  OAI21X1 U20062 ( .A(n27094), .B(n29219), .C(n23832), .Y(n30176) );
  AOI22X1 U20063 ( .A(n30174), .B(n29217), .C(net64168), .D(n30176), .Y(n30177) );
  AOI22X1 U20064 ( .A(n30954), .B(n29320), .C(n29441), .D(n32270), .Y(n30184)
         );
  AOI21X1 U20065 ( .A(n23325), .B(n34498), .C(n30180), .Y(n30181) );
  OAI21X1 U20066 ( .A(n27092), .B(n29219), .C(n23833), .Y(n30182) );
  AOI22X1 U20067 ( .A(n30180), .B(n29217), .C(net64168), .D(n30182), .Y(n30183) );
  NAND3X1 U20068 ( .A(data_in[4]), .B(n30371), .C(n30234), .Y(n30185) );
  NAND3X1 U20069 ( .A(n21186), .B(n30186), .C(n26271), .Y(n30187) );
  AOI22X1 U20070 ( .A(n30975), .B(n29320), .C(n29441), .D(n32275), .Y(n30194)
         );
  NAND3X1 U20071 ( .A(n29461), .B(n33996), .C(n25451), .Y(n30188) );
  NAND3X1 U20072 ( .A(net53623), .B(n29443), .C(net104479), .Y(n30189) );
  AOI21X1 U20073 ( .A(n23328), .B(n34498), .C(n30190), .Y(n30191) );
  OAI21X1 U20074 ( .A(n25358), .B(n29219), .C(n23834), .Y(n30192) );
  AOI22X1 U20075 ( .A(n30190), .B(n29217), .C(net64168), .D(n30192), .Y(n30193) );
  AOI22X1 U20076 ( .A(n31001), .B(n29320), .C(n29440), .D(n23329), .Y(n30199)
         );
  AOI21X1 U20077 ( .A(n23330), .B(n34498), .C(n30195), .Y(n30196) );
  OAI21X1 U20078 ( .A(n26873), .B(n29219), .C(n23835), .Y(n30197) );
  AOI22X1 U20079 ( .A(n30195), .B(n29217), .C(net64168), .D(n30197), .Y(n30198) );
  AOI22X1 U20080 ( .A(n31011), .B(n29320), .C(n29440), .D(n32283), .Y(n30204)
         );
  AOI21X1 U20081 ( .A(n23333), .B(n34498), .C(n30200), .Y(n30201) );
  OAI21X1 U20082 ( .A(n25359), .B(n29219), .C(n23836), .Y(n30202) );
  AOI22X1 U20083 ( .A(n30200), .B(n29217), .C(net64168), .D(n30202), .Y(n30203) );
  AOI22X1 U20084 ( .A(n31038), .B(n29320), .C(n29441), .D(n23334), .Y(n30209)
         );
  AOI21X1 U20085 ( .A(n23335), .B(n34498), .C(n30205), .Y(n30206) );
  OAI21X1 U20086 ( .A(n26759), .B(n29219), .C(n23837), .Y(n30207) );
  AOI22X1 U20087 ( .A(n30205), .B(n29217), .C(net64168), .D(n30207), .Y(n30208) );
  AOI22X1 U20088 ( .A(n31049), .B(n29320), .C(n29440), .D(n32291), .Y(n30214)
         );
  AOI21X1 U20089 ( .A(n23337), .B(n34498), .C(n30210), .Y(n30211) );
  OAI21X1 U20090 ( .A(n25360), .B(n29219), .C(n23838), .Y(n30212) );
  AOI22X1 U20091 ( .A(n30210), .B(n29217), .C(net64168), .D(n30212), .Y(n30213) );
  AOI22X1 U20092 ( .A(n31076), .B(n29320), .C(n29441), .D(n23338), .Y(n30219)
         );
  AOI21X1 U20093 ( .A(n23339), .B(n34498), .C(n30215), .Y(n30216) );
  OAI21X1 U20094 ( .A(n27111), .B(n29219), .C(n23839), .Y(n30217) );
  AOI22X1 U20095 ( .A(n30215), .B(n29217), .C(net64168), .D(n30217), .Y(n30218) );
  AOI22X1 U20096 ( .A(n31089), .B(n29320), .C(n29441), .D(n32299), .Y(n30224)
         );
  AOI21X1 U20097 ( .A(n23341), .B(n34498), .C(n30220), .Y(n30221) );
  OAI21X1 U20098 ( .A(n25361), .B(n29219), .C(n23840), .Y(n30222) );
  AOI22X1 U20099 ( .A(n30220), .B(n29217), .C(net64168), .D(n30222), .Y(n30223) );
  AOI22X1 U20100 ( .A(n31116), .B(n29320), .C(n29440), .D(n23342), .Y(n30233)
         );
  AOI21X1 U20101 ( .A(n23343), .B(n34498), .C(n30229), .Y(n30230) );
  OAI21X1 U20102 ( .A(n27014), .B(n29219), .C(n23841), .Y(n30231) );
  AOI22X1 U20103 ( .A(n30229), .B(n29217), .C(net64168), .D(n30231), .Y(n30232) );
  NAND3X1 U20104 ( .A(data_in[4]), .B(data_in[3]), .C(n30234), .Y(n30235) );
  AOI22X1 U20105 ( .A(n31129), .B(n29320), .C(n29440), .D(n32307), .Y(n30242)
         );
  NAND3X1 U20106 ( .A(n25451), .B(n33996), .C(n28606), .Y(n30236) );
  NAND3X1 U20107 ( .A(net53623), .B(net104479), .C(n28220), .Y(n30237) );
  AOI21X1 U20108 ( .A(n23345), .B(n34498), .C(n30238), .Y(n30239) );
  OAI21X1 U20109 ( .A(n25362), .B(n29219), .C(n23842), .Y(n30240) );
  AOI22X1 U20110 ( .A(n30238), .B(n29217), .C(net64168), .D(n30240), .Y(n30241) );
  AOI22X1 U20111 ( .A(n31156), .B(n29320), .C(n29441), .D(n23346), .Y(n30247)
         );
  AOI21X1 U20112 ( .A(n23456), .B(n34498), .C(n30243), .Y(n30244) );
  OAI21X1 U20113 ( .A(n26814), .B(n29219), .C(n23843), .Y(n30245) );
  AOI22X1 U20114 ( .A(n30243), .B(n29217), .C(net64168), .D(n30245), .Y(n30246) );
  AOI22X1 U20115 ( .A(n31167), .B(n29320), .C(n29441), .D(n32315), .Y(n30252)
         );
  AOI21X1 U20116 ( .A(n23348), .B(n34498), .C(n30248), .Y(n30249) );
  OAI21X1 U20117 ( .A(n25342), .B(n29219), .C(n23844), .Y(n30250) );
  AOI22X1 U20118 ( .A(n30248), .B(n29217), .C(net64168), .D(n30250), .Y(n30251) );
  AOI22X1 U20119 ( .A(n31193), .B(n29320), .C(n29440), .D(n23349), .Y(n30257)
         );
  AOI21X1 U20120 ( .A(n23350), .B(n34498), .C(n30253), .Y(n30254) );
  OAI21X1 U20121 ( .A(n27108), .B(n29219), .C(n23845), .Y(n30255) );
  AOI22X1 U20122 ( .A(n30253), .B(n29217), .C(net64168), .D(n30255), .Y(n30256) );
  AOI22X1 U20123 ( .A(n31206), .B(n29320), .C(n29441), .D(n32323), .Y(n30262)
         );
  AOI21X1 U20124 ( .A(n23352), .B(n34498), .C(n30258), .Y(n30259) );
  OAI21X1 U20125 ( .A(n25363), .B(n29219), .C(n23846), .Y(n30260) );
  AOI22X1 U20126 ( .A(n30258), .B(n29217), .C(net64168), .D(n30260), .Y(n30261) );
  AOI22X1 U20127 ( .A(n31233), .B(n29320), .C(n29440), .D(n23353), .Y(n30267)
         );
  AOI21X1 U20128 ( .A(n23354), .B(n34498), .C(n30263), .Y(n30264) );
  OAI21X1 U20129 ( .A(n27011), .B(n29219), .C(n23847), .Y(n30265) );
  AOI22X1 U20130 ( .A(n30263), .B(n29217), .C(net64168), .D(n30265), .Y(n30266) );
  AOI22X1 U20131 ( .A(n31246), .B(n29320), .C(n29441), .D(n32331), .Y(n30271)
         );
  AOI21X1 U20132 ( .A(n23356), .B(n34498), .C(n34606), .Y(n30268) );
  OAI21X1 U20133 ( .A(n25364), .B(n29219), .C(n23848), .Y(n30269) );
  AOI22X1 U20134 ( .A(n34606), .B(n29217), .C(net64168), .D(n30269), .Y(n30270) );
  AOI22X1 U20135 ( .A(n31273), .B(n29320), .C(n29440), .D(n21169), .Y(n30279)
         );
  AOI21X1 U20136 ( .A(n23357), .B(n34498), .C(n30275), .Y(n30276) );
  OAI21X1 U20137 ( .A(n26946), .B(n29219), .C(n23849), .Y(n30277) );
  AOI22X1 U20138 ( .A(n30275), .B(n29217), .C(net64168), .D(n30277), .Y(n30278) );
  NAND3X1 U20139 ( .A(data_in[5]), .B(n30371), .C(n30327), .Y(n30280) );
  AOI22X1 U20140 ( .A(n32045), .B(n29320), .C(n29440), .D(n32339), .Y(n30288)
         );
  NAND3X1 U20141 ( .A(n29461), .B(n33995), .C(n27210), .Y(n30282) );
  NAND3X1 U20142 ( .A(net53601), .B(n29443), .C(net124030), .Y(n30283) );
  AOI21X1 U20143 ( .A(n23359), .B(n34498), .C(n30284), .Y(n30285) );
  OAI21X1 U20144 ( .A(n25365), .B(n29219), .C(n23850), .Y(n30286) );
  AOI22X1 U20145 ( .A(n30284), .B(n29217), .C(net64168), .D(n30286), .Y(n30287) );
  AOI22X1 U20146 ( .A(n31303), .B(n29320), .C(n29441), .D(n32343), .Y(n30293)
         );
  AOI21X1 U20147 ( .A(n23361), .B(n34498), .C(n30289), .Y(n30290) );
  OAI21X1 U20148 ( .A(n25366), .B(n29219), .C(n23851), .Y(n30291) );
  AOI22X1 U20149 ( .A(n30289), .B(n29217), .C(net64168), .D(n30291), .Y(n30292) );
  AOI22X1 U20150 ( .A(n32053), .B(n29320), .C(n29441), .D(n32347), .Y(n30298)
         );
  AOI21X1 U20151 ( .A(n23363), .B(n34498), .C(n30294), .Y(n30295) );
  OAI21X1 U20152 ( .A(n25367), .B(n29219), .C(n23852), .Y(n30296) );
  AOI22X1 U20153 ( .A(n30294), .B(n29217), .C(net64168), .D(n30296), .Y(n30297) );
  AOI22X1 U20154 ( .A(n31340), .B(n29320), .C(n29440), .D(n32351), .Y(n30303)
         );
  AOI21X1 U20155 ( .A(n23366), .B(n34498), .C(n30299), .Y(n30300) );
  OAI21X1 U20156 ( .A(n25368), .B(n29219), .C(n23853), .Y(n30301) );
  AOI22X1 U20157 ( .A(n30299), .B(n29217), .C(net64168), .D(n30301), .Y(n30302) );
  AOI22X1 U20158 ( .A(n32060), .B(n29320), .C(n29440), .D(n32355), .Y(n30308)
         );
  AOI21X1 U20159 ( .A(n23368), .B(n34498), .C(n30304), .Y(n30305) );
  OAI21X1 U20160 ( .A(n25369), .B(n29219), .C(n23854), .Y(n30306) );
  AOI22X1 U20161 ( .A(n30304), .B(n29217), .C(net64168), .D(n30306), .Y(n30307) );
  AOI22X1 U20162 ( .A(n31380), .B(n29320), .C(n29440), .D(n32359), .Y(n30313)
         );
  AOI21X1 U20163 ( .A(n23370), .B(n34498), .C(n30309), .Y(n30310) );
  OAI21X1 U20164 ( .A(n25370), .B(n29219), .C(n23855), .Y(n30311) );
  AOI22X1 U20165 ( .A(n30309), .B(n29217), .C(net64168), .D(n30311), .Y(n30312) );
  AOI22X1 U20166 ( .A(n32068), .B(n29320), .C(n29440), .D(n32363), .Y(n30318)
         );
  AOI21X1 U20167 ( .A(n23372), .B(n34498), .C(n30314), .Y(n30315) );
  OAI21X1 U20168 ( .A(n25371), .B(n29219), .C(n23856), .Y(n30316) );
  AOI22X1 U20169 ( .A(n30314), .B(n29217), .C(net64168), .D(n30316), .Y(n30317) );
  AOI22X1 U20170 ( .A(n31421), .B(n29320), .C(n29440), .D(n32367), .Y(n30326)
         );
  AOI21X1 U20171 ( .A(n23374), .B(n34498), .C(n30322), .Y(n30323) );
  OAI21X1 U20172 ( .A(n25372), .B(n29219), .C(n23857), .Y(n30324) );
  AOI22X1 U20173 ( .A(n30322), .B(n29217), .C(net64168), .D(n30324), .Y(n30325) );
  AOI22X1 U20174 ( .A(n32076), .B(n29320), .C(n29440), .D(n32371), .Y(n30334)
         );
  NAND3X1 U20175 ( .A(n27210), .B(n33995), .C(n28606), .Y(n30328) );
  NAND3X1 U20176 ( .A(net53601), .B(net124030), .C(n28220), .Y(n30329) );
  AOI21X1 U20177 ( .A(n23376), .B(n34498), .C(n30330), .Y(n30331) );
  OAI21X1 U20178 ( .A(n25373), .B(n29219), .C(n23858), .Y(n30332) );
  AOI22X1 U20179 ( .A(n30330), .B(n29217), .C(net64168), .D(n30332), .Y(n30333) );
  AOI22X1 U20180 ( .A(n31460), .B(n29320), .C(n29440), .D(n32375), .Y(n30339)
         );
  AOI21X1 U20181 ( .A(n23378), .B(n34498), .C(n30335), .Y(n30336) );
  OAI21X1 U20182 ( .A(n25374), .B(n29219), .C(n23859), .Y(n30337) );
  AOI22X1 U20183 ( .A(n30335), .B(n29217), .C(net64168), .D(n30337), .Y(n30338) );
  AOI22X1 U20184 ( .A(n32084), .B(n29320), .C(n29440), .D(n32379), .Y(n30344)
         );
  AOI21X1 U20185 ( .A(n23380), .B(n34498), .C(n30340), .Y(n30341) );
  OAI21X1 U20186 ( .A(n25375), .B(n29219), .C(n23860), .Y(n30342) );
  AOI22X1 U20187 ( .A(n30340), .B(n29217), .C(net64168), .D(n30342), .Y(n30343) );
  AOI22X1 U20188 ( .A(n31499), .B(n29320), .C(n29440), .D(n32383), .Y(n30348)
         );
  AOI21X1 U20189 ( .A(n23383), .B(n34498), .C(n34609), .Y(n30345) );
  OAI21X1 U20190 ( .A(n25376), .B(n29219), .C(n23861), .Y(n30346) );
  AOI22X1 U20191 ( .A(n34609), .B(n29217), .C(net64168), .D(n30346), .Y(n30347) );
  AOI22X1 U20192 ( .A(n32091), .B(n29320), .C(n29440), .D(n32387), .Y(n30353)
         );
  AOI21X1 U20193 ( .A(n23385), .B(n34498), .C(n30349), .Y(n30350) );
  OAI21X1 U20194 ( .A(n25377), .B(n29219), .C(n23862), .Y(n30351) );
  AOI22X1 U20195 ( .A(n30349), .B(n29217), .C(net64168), .D(n30351), .Y(n30352) );
  AOI22X1 U20196 ( .A(n31537), .B(n29320), .C(n29440), .D(n32391), .Y(n30358)
         );
  AOI21X1 U20197 ( .A(n23387), .B(n34498), .C(n30354), .Y(n30355) );
  OAI21X1 U20198 ( .A(n25378), .B(n29219), .C(n23863), .Y(n30356) );
  AOI22X1 U20199 ( .A(n30354), .B(n29217), .C(net64168), .D(n30356), .Y(n30357) );
  AOI22X1 U20200 ( .A(n32100), .B(n29320), .C(n29440), .D(n32395), .Y(n30363)
         );
  AOI21X1 U20201 ( .A(n23389), .B(n34498), .C(n30359), .Y(n30360) );
  OAI21X1 U20202 ( .A(n25379), .B(n29219), .C(n23864), .Y(n30361) );
  AOI22X1 U20203 ( .A(n30359), .B(n29217), .C(net64168), .D(n30361), .Y(n30362) );
  AOI22X1 U20204 ( .A(n31578), .B(n29320), .C(n29440), .D(n32399), .Y(n30370)
         );
  AOI21X1 U20205 ( .A(n23391), .B(n34498), .C(n30366), .Y(n30367) );
  OAI21X1 U20206 ( .A(n25380), .B(n29219), .C(n23865), .Y(n30368) );
  AOI22X1 U20207 ( .A(n30366), .B(n29217), .C(net64168), .D(n30368), .Y(n30369) );
  NAND3X1 U20208 ( .A(data_in[5]), .B(data_in[4]), .C(n30371), .Y(n30372) );
  AOI22X1 U20209 ( .A(n31598), .B(n29320), .C(n29441), .D(n32403), .Y(n30379)
         );
  NAND3X1 U20210 ( .A(n27211), .B(n29461), .C(n25451), .Y(n30373) );
  NAND3X1 U20211 ( .A(n29443), .B(net124030), .C(net104479), .Y(n30374) );
  AOI21X1 U20212 ( .A(n23393), .B(n34498), .C(n30375), .Y(n30376) );
  OAI21X1 U20213 ( .A(n25381), .B(n29219), .C(n23866), .Y(n30377) );
  AOI22X1 U20214 ( .A(n30375), .B(n29217), .C(net64168), .D(n30377), .Y(n30378) );
  AOI22X1 U20215 ( .A(n31624), .B(n29320), .C(n29441), .D(n23394), .Y(n30384)
         );
  AOI21X1 U20216 ( .A(n23395), .B(n34498), .C(n30380), .Y(n30381) );
  OAI21X1 U20217 ( .A(n25383), .B(n29219), .C(n23867), .Y(n30382) );
  AOI22X1 U20218 ( .A(n30380), .B(n29217), .C(net64168), .D(n30382), .Y(n30383) );
  AOI22X1 U20219 ( .A(n31635), .B(n29320), .C(n29441), .D(n32411), .Y(n30388)
         );
  AOI21X1 U20220 ( .A(n23397), .B(n34498), .C(n34599), .Y(n30385) );
  OAI21X1 U20221 ( .A(n25384), .B(n29219), .C(n23868), .Y(n30386) );
  AOI22X1 U20222 ( .A(n34599), .B(n29217), .C(net64168), .D(n30386), .Y(n30387) );
  AOI22X1 U20223 ( .A(n31660), .B(n29320), .C(n29441), .D(n23398), .Y(n30393)
         );
  AOI21X1 U20224 ( .A(n23399), .B(n34498), .C(n30389), .Y(n30390) );
  OAI21X1 U20225 ( .A(n27009), .B(n29219), .C(n23869), .Y(n30391) );
  AOI22X1 U20226 ( .A(n30389), .B(n29217), .C(net64168), .D(n30391), .Y(n30392) );
  AOI22X1 U20227 ( .A(n31672), .B(n29320), .C(n29441), .D(n32419), .Y(n30398)
         );
  AOI21X1 U20228 ( .A(n23401), .B(n34498), .C(n30394), .Y(n30395) );
  OAI21X1 U20229 ( .A(n25385), .B(n29219), .C(n23870), .Y(n30396) );
  AOI22X1 U20230 ( .A(n30394), .B(n29217), .C(net64168), .D(n30396), .Y(n30397) );
  AOI22X1 U20231 ( .A(n31698), .B(n29320), .C(n29441), .D(n23402), .Y(n30403)
         );
  AOI21X1 U20232 ( .A(n23403), .B(n34498), .C(n30399), .Y(n30400) );
  OAI21X1 U20233 ( .A(n26944), .B(n29219), .C(n23871), .Y(n30401) );
  AOI22X1 U20234 ( .A(n30399), .B(n29217), .C(net64168), .D(n30401), .Y(n30402) );
  AOI22X1 U20235 ( .A(n31711), .B(n29320), .C(n29441), .D(n32427), .Y(n30408)
         );
  AOI21X1 U20236 ( .A(n23405), .B(n34498), .C(n30404), .Y(n30405) );
  OAI21X1 U20237 ( .A(n25386), .B(n29219), .C(n23872), .Y(n30406) );
  AOI22X1 U20238 ( .A(n30404), .B(n29217), .C(net64168), .D(n30406), .Y(n30407) );
  AOI22X1 U20239 ( .A(n31738), .B(n29320), .C(n29441), .D(n23406), .Y(n30417)
         );
  AOI21X1 U20240 ( .A(n23408), .B(n34498), .C(n30413), .Y(n30414) );
  OAI21X1 U20241 ( .A(n25387), .B(n29219), .C(n23873), .Y(n30415) );
  AOI22X1 U20242 ( .A(n30413), .B(n29217), .C(net64168), .D(n30415), .Y(n30416) );
  AOI22X1 U20243 ( .A(n31749), .B(n29320), .C(n29441), .D(n32434), .Y(n30425)
         );
  NAND3X1 U20244 ( .A(n25451), .B(n27210), .C(n28606), .Y(n30419) );
  NAND3X1 U20245 ( .A(net104479), .B(net124030), .C(n28220), .Y(n30420) );
  AOI21X1 U20246 ( .A(n23410), .B(n34498), .C(n30421), .Y(n30422) );
  OAI21X1 U20247 ( .A(n25388), .B(n29219), .C(n23874), .Y(n30423) );
  AOI22X1 U20248 ( .A(n30421), .B(n29217), .C(net64168), .D(n30423), .Y(n30424) );
  AOI22X1 U20249 ( .A(n31776), .B(n29320), .C(n29441), .D(n23411), .Y(n30431)
         );
  AOI21X1 U20250 ( .A(n23412), .B(n34498), .C(n30427), .Y(n30428) );
  OAI21X1 U20251 ( .A(n27105), .B(n29219), .C(n23875), .Y(n30429) );
  AOI22X1 U20252 ( .A(n30427), .B(n29217), .C(net64168), .D(n30429), .Y(n30430) );
  AOI22X1 U20253 ( .A(n31789), .B(n29320), .C(n29441), .D(n32442), .Y(n30439)
         );
  AOI21X1 U20254 ( .A(n23414), .B(n34498), .C(n30435), .Y(n30436) );
  OAI21X1 U20255 ( .A(n25389), .B(n29219), .C(n23876), .Y(n30437) );
  AOI22X1 U20256 ( .A(n30435), .B(n29217), .C(net64168), .D(n30437), .Y(n30438) );
  AOI22X1 U20257 ( .A(n31815), .B(n29320), .C(n29441), .D(n23415), .Y(n30448)
         );
  AOI21X1 U20258 ( .A(n23416), .B(n34498), .C(n30444), .Y(n30445) );
  OAI21X1 U20259 ( .A(n26943), .B(n29219), .C(n23877), .Y(n30446) );
  AOI22X1 U20260 ( .A(n30444), .B(n29217), .C(net64168), .D(n30446), .Y(n30447) );
  AOI22X1 U20261 ( .A(n31828), .B(n29320), .C(n29441), .D(n32450), .Y(n30456)
         );
  AOI21X1 U20262 ( .A(n23418), .B(n34498), .C(n30452), .Y(n30453) );
  OAI21X1 U20263 ( .A(n25390), .B(n29219), .C(n23878), .Y(n30454) );
  AOI22X1 U20264 ( .A(n30452), .B(n29217), .C(net64168), .D(n30454), .Y(n30455) );
  AOI22X1 U20265 ( .A(n31855), .B(n29320), .C(n29440), .D(n23419), .Y(n30463)
         );
  AOI21X1 U20266 ( .A(n23421), .B(n34498), .C(n34602), .Y(n30460) );
  OAI21X1 U20267 ( .A(n25391), .B(n29219), .C(n23879), .Y(n30461) );
  AOI22X1 U20268 ( .A(n34602), .B(n29217), .C(net64168), .D(n30461), .Y(n30462) );
  AOI22X1 U20269 ( .A(n31867), .B(n29320), .C(n29441), .D(n32457), .Y(n30470)
         );
  AOI21X1 U20270 ( .A(n23423), .B(n34498), .C(n30466), .Y(n30467) );
  OAI21X1 U20271 ( .A(n25392), .B(n29219), .C(n23880), .Y(n30468) );
  AOI22X1 U20272 ( .A(n30466), .B(n29217), .C(net64168), .D(n30468), .Y(n30469) );
  OAI21X1 U20273 ( .A(n29219), .B(n25434), .C(n24963), .Y(n30477) );
  OAI21X1 U20274 ( .A(n24280), .B(n30477), .C(net64168), .Y(n30479) );
  OAI21X1 U20275 ( .A(n27062), .B(n27179), .C(n23890), .Y(n30483) );
  INVX2 U20276 ( .A(n14097), .Y(n30487) );
  NOR2X1 U20277 ( .A(n24983), .B(n30487), .Y(n14351) );
  INVX2 U20278 ( .A(n14373), .Y(n30616) );
  NAND2X1 U20279 ( .A(n30021), .B(n30616), .Y(n30488) );
  NAND2X1 U20280 ( .A(n29352), .B(n30616), .Y(n32190) );
  AOI22X1 U20281 ( .A(n29337), .B(n24928), .C(n29334), .D(n30489), .Y(n30493)
         );
  NAND2X1 U20282 ( .A(n30038), .B(n30616), .Y(n30490) );
  AOI22X1 U20283 ( .A(n29340), .B(n33875), .C(n25083), .D(n30616), .Y(n30492)
         );
  NAND2X1 U20284 ( .A(n30493), .B(n30492), .Y(n15851) );
  AOI22X1 U20285 ( .A(n29336), .B(n27079), .C(n29334), .D(n30494), .Y(n30498)
         );
  AOI22X1 U20286 ( .A(n29340), .B(n33852), .C(n26980), .D(n30616), .Y(n30497)
         );
  NAND2X1 U20287 ( .A(n30498), .B(n30497), .Y(n15830) );
  AOI22X1 U20288 ( .A(n29336), .B(n23614), .C(n29334), .D(n30499), .Y(n30502)
         );
  AOI22X1 U20289 ( .A(n29340), .B(n33829), .C(n26594), .D(n30616), .Y(n30501)
         );
  NAND2X1 U20290 ( .A(n30502), .B(n30501), .Y(n15809) );
  AOI22X1 U20291 ( .A(n29336), .B(n26997), .C(n29333), .D(n30503), .Y(n30507)
         );
  AOI22X1 U20292 ( .A(n29340), .B(n33806), .C(n26619), .D(n30616), .Y(n30506)
         );
  NAND2X1 U20293 ( .A(n30507), .B(n30506), .Y(n15788) );
  AOI22X1 U20294 ( .A(n29336), .B(n27174), .C(n29333), .D(n30508), .Y(n30512)
         );
  AOI22X1 U20295 ( .A(n29340), .B(n33784), .C(n26645), .D(n30616), .Y(n30511)
         );
  NAND2X1 U20296 ( .A(n30512), .B(n30511), .Y(n15767) );
  AOI22X1 U20297 ( .A(n29336), .B(n22943), .C(n29333), .D(n30513), .Y(n30517)
         );
  AOI22X1 U20298 ( .A(n29340), .B(n33762), .C(n26677), .D(n30616), .Y(n30516)
         );
  NAND2X1 U20299 ( .A(n30517), .B(n30516), .Y(n15746) );
  AOI22X1 U20300 ( .A(n29336), .B(n22944), .C(n29333), .D(n30518), .Y(n30522)
         );
  AOI22X1 U20301 ( .A(n29340), .B(n26077), .C(n26709), .D(n30616), .Y(n30521)
         );
  NAND2X1 U20302 ( .A(n30522), .B(n30521), .Y(n15724) );
  AOI22X1 U20303 ( .A(n29336), .B(n24929), .C(n29333), .D(n30523), .Y(n30526)
         );
  AOI22X1 U20304 ( .A(n29340), .B(n33718), .C(n26796), .D(n30616), .Y(n30525)
         );
  NAND2X1 U20305 ( .A(n30526), .B(n30525), .Y(n15702) );
  AOI22X1 U20306 ( .A(n29336), .B(n24930), .C(n29333), .D(n30527), .Y(n30530)
         );
  AOI22X1 U20307 ( .A(n29340), .B(n33696), .C(n26751), .D(n30616), .Y(n30529)
         );
  NAND2X1 U20308 ( .A(n30530), .B(n30529), .Y(n15681) );
  AOI22X1 U20309 ( .A(n29336), .B(n24931), .C(n29333), .D(n30531), .Y(n30534)
         );
  AOI22X1 U20310 ( .A(n29340), .B(n33661), .C(n26850), .D(n30616), .Y(n30533)
         );
  NAND2X1 U20311 ( .A(n30534), .B(n30533), .Y(n15660) );
  AOI22X1 U20312 ( .A(n29336), .B(n22945), .C(n29333), .D(n30535), .Y(n30539)
         );
  AOI22X1 U20313 ( .A(n29340), .B(n33653), .C(n25084), .D(n30616), .Y(n30538)
         );
  NAND2X1 U20314 ( .A(n30539), .B(n30538), .Y(n15639) );
  AOI22X1 U20315 ( .A(n29336), .B(n22946), .C(n29333), .D(n30540), .Y(n30544)
         );
  AOI22X1 U20316 ( .A(n29341), .B(n21232), .C(n26913), .D(n30616), .Y(n30543)
         );
  NAND2X1 U20317 ( .A(n30544), .B(n30543), .Y(n15618) );
  AOI22X1 U20318 ( .A(n29337), .B(n22949), .C(n29333), .D(n30545), .Y(n30549)
         );
  AOI22X1 U20319 ( .A(n29340), .B(n33609), .C(n27161), .D(n30616), .Y(n30548)
         );
  NAND2X1 U20320 ( .A(n30549), .B(n30548), .Y(n15597) );
  OAI21X1 U20321 ( .A(n30062), .B(n25432), .C(n25106), .Y(n30552) );
  AOI22X1 U20322 ( .A(n30552), .B(n30616), .C(n29336), .D(n26521), .Y(n30553)
         );
  OAI21X1 U20323 ( .A(n30554), .B(n32190), .C(n30553), .Y(n15580) );
  OAI21X1 U20324 ( .A(n33531), .B(n25082), .C(n29341), .Y(n30560) );
  NAND2X1 U20325 ( .A(n30556), .B(n30616), .Y(n33561) );
  AOI22X1 U20326 ( .A(n29337), .B(n22951), .C(n29333), .D(n30557), .Y(n30559)
         );
  NAND3X1 U20327 ( .A(n30560), .B(n33561), .C(n30559), .Y(n15529) );
  OAI21X1 U20328 ( .A(n33508), .B(n25134), .C(n29341), .Y(n30564) );
  AOI22X1 U20329 ( .A(n29337), .B(n23633), .C(n29333), .D(n30562), .Y(n30563)
         );
  NAND3X1 U20330 ( .A(n30564), .B(n33561), .C(n30563), .Y(n15508) );
  OAI21X1 U20331 ( .A(n33485), .B(n25135), .C(n29341), .Y(n30569) );
  AOI22X1 U20332 ( .A(n29337), .B(n22952), .C(n29332), .D(n30566), .Y(n30568)
         );
  NAND3X1 U20333 ( .A(n30569), .B(n33561), .C(n30568), .Y(n15486) );
  OAI21X1 U20334 ( .A(n33462), .B(n25136), .C(n29341), .Y(n30574) );
  AOI22X1 U20335 ( .A(n29337), .B(n22953), .C(n29332), .D(n30571), .Y(n30573)
         );
  NAND3X1 U20336 ( .A(n30574), .B(n33561), .C(n30573), .Y(n15464) );
  OAI21X1 U20337 ( .A(n25774), .B(n25137), .C(n29341), .Y(n30579) );
  AOI22X1 U20338 ( .A(n29337), .B(n22954), .C(n29332), .D(n30576), .Y(n30578)
         );
  NAND3X1 U20339 ( .A(n30579), .B(n33561), .C(n30578), .Y(n15442) );
  OAI21X1 U20340 ( .A(n33417), .B(n25138), .C(n29341), .Y(n30584) );
  AOI22X1 U20341 ( .A(n29337), .B(n22955), .C(n29332), .D(n30581), .Y(n30583)
         );
  NAND3X1 U20342 ( .A(n30584), .B(n33561), .C(n30583), .Y(n15420) );
  OAI21X1 U20343 ( .A(n25657), .B(n25139), .C(n29341), .Y(n30589) );
  AOI22X1 U20344 ( .A(n29337), .B(n22956), .C(n29332), .D(n30586), .Y(n30588)
         );
  NAND3X1 U20345 ( .A(n30589), .B(n33561), .C(n30588), .Y(n15397) );
  OAI21X1 U20346 ( .A(n25680), .B(n25140), .C(n29341), .Y(n30594) );
  AOI22X1 U20347 ( .A(n29337), .B(n22957), .C(n29332), .D(n30591), .Y(n30593)
         );
  NAND3X1 U20348 ( .A(n30594), .B(n33561), .C(n30593), .Y(n15373) );
  OAI21X1 U20349 ( .A(n33326), .B(n25141), .C(n29341), .Y(n30599) );
  AOI22X1 U20350 ( .A(n29337), .B(n22958), .C(n29332), .D(n30596), .Y(n30598)
         );
  NAND3X1 U20351 ( .A(n30599), .B(n33561), .C(n30598), .Y(n15348) );
  OAI21X1 U20352 ( .A(n33295), .B(n25142), .C(n29341), .Y(n30604) );
  AOI22X1 U20353 ( .A(n29337), .B(n22959), .C(n29332), .D(n30601), .Y(n30603)
         );
  NAND3X1 U20354 ( .A(n30604), .B(n33561), .C(n30603), .Y(n15325) );
  OAI21X1 U20355 ( .A(n25658), .B(n25143), .C(n29341), .Y(n30609) );
  AOI22X1 U20356 ( .A(n29337), .B(n22960), .C(n29332), .D(n30606), .Y(n30608)
         );
  NAND3X1 U20357 ( .A(n30609), .B(n33561), .C(n30608), .Y(n15302) );
  OAI21X1 U20358 ( .A(n33234), .B(n25144), .C(n29341), .Y(n30614) );
  AOI22X1 U20359 ( .A(n29338), .B(n22961), .C(n29332), .D(n30611), .Y(n30613)
         );
  NAND3X1 U20360 ( .A(n30614), .B(n33561), .C(n30613), .Y(n15279) );
  NAND2X1 U20361 ( .A(n29341), .B(n25118), .Y(n30620) );
  NAND2X1 U20362 ( .A(n30617), .B(n30616), .Y(n30624) );
  AOI22X1 U20363 ( .A(n29338), .B(n25006), .C(n29332), .D(n30618), .Y(n30619)
         );
  NAND3X1 U20364 ( .A(n30620), .B(n30624), .C(n30619), .Y(n15256) );
  OAI21X1 U20365 ( .A(n32764), .B(n34342), .C(n29341), .Y(n30621) );
  OAI21X1 U20366 ( .A(n30622), .B(n32190), .C(n30621), .Y(n30623) );
  OAI21X1 U20367 ( .A(n34342), .B(n34222), .C(n29338), .Y(n30625) );
  NAND3X1 U20368 ( .A(n30628), .B(n30625), .C(n30624), .Y(n15235) );
  AOI22X1 U20369 ( .A(n29338), .B(n25068), .C(n29340), .D(n23457), .Y(n30627)
         );
  NAND3X1 U20370 ( .A(n30628), .B(n33561), .C(n30627), .Y(n15226) );
  OAI21X1 U20371 ( .A(n29191), .B(n34555), .C(net64168), .Y(n30629) );
  AOI21X1 U20372 ( .A(n24269), .B(n27196), .C(n21408), .Y(n31890) );
  AOI22X1 U20373 ( .A(n26315), .B(n23311), .C(n26020), .D(n25715), .Y(n30649)
         );
  OAI21X1 U20374 ( .A(n25846), .B(n21072), .C(n23443), .Y(n30639) );
  AOI21X1 U20375 ( .A(n29269), .B(n25357), .C(n20839), .Y(n30640) );
  OAI21X1 U20376 ( .A(n23311), .B(n29260), .C(n21926), .Y(n30641) );
  NAND3X1 U20377 ( .A(n30644), .B(n30643), .C(n30642), .Y(n31913) );
  OAI21X1 U20378 ( .A(n25715), .B(n29254), .C(n26331), .Y(n30645) );
  AOI21X1 U20379 ( .A(n26465), .B(n23310), .C(n22150), .Y(n30647) );
  NAND3X1 U20380 ( .A(n24047), .B(n23458), .C(n22795), .Y(n22055) );
  OAI21X1 U20381 ( .A(locTrig[3]), .B(n21170), .C(n30636), .Y(n31901) );
  AOI22X1 U20382 ( .A(n20819), .B(n23310), .C(n25536), .D(n23311), .Y(n30662)
         );
  AOI21X1 U20383 ( .A(n24270), .B(n30653), .C(n21408), .Y(n31899) );
  OAI21X1 U20384 ( .A(n30655), .B(n29237), .C(n22998), .Y(n30659) );
  NOR3X1 U20385 ( .A(n30659), .B(n29285), .C(n30664), .Y(n30660) );
  NAND3X1 U20386 ( .A(n30660), .B(n24446), .C(n22735), .Y(n22054) );
  OAI21X1 U20387 ( .A(n27181), .B(n30663), .C(n24936), .Y(n31885) );
  AOI21X1 U20388 ( .A(n25854), .B(n25715), .C(n30658), .Y(n30669) );
  OAI21X1 U20389 ( .A(n23279), .B(net149842), .C(n30631), .Y(n30665) );
  OAI21X1 U20390 ( .A(n30655), .B(n29319), .C(n29210), .Y(n30666) );
  AOI21X1 U20391 ( .A(n25799), .B(n23311), .C(n30666), .Y(n30667) );
  NAND3X1 U20392 ( .A(n25224), .B(n24848), .C(n22727), .Y(n22053) );
  AOI22X1 U20393 ( .A(n26309), .B(n23312), .C(n26040), .D(n32199), .Y(n30677)
         );
  AOI21X1 U20394 ( .A(n29269), .B(n26935), .C(n26293), .Y(n30671) );
  OAI21X1 U20395 ( .A(n23312), .B(n29260), .C(n21927), .Y(n30672) );
  OAI21X1 U20396 ( .A(n32199), .B(n29254), .C(n26324), .Y(n30673) );
  AOI21X1 U20397 ( .A(n26462), .B(n32200), .C(n22154), .Y(n30675) );
  AOI22X1 U20398 ( .A(n29197), .B(n32200), .C(n25549), .D(n23312), .Y(n30682)
         );
  OAI21X1 U20399 ( .A(n30683), .B(n29237), .C(n23189), .Y(n30679) );
  NOR3X1 U20400 ( .A(n30679), .B(n29283), .C(n30678), .Y(n30680) );
  NAND3X1 U20401 ( .A(n24447), .B(n30680), .C(n22286), .Y(n22060) );
  AOI21X1 U20402 ( .A(n29315), .B(n27166), .C(n29278), .Y(n30693) );
  OAI21X1 U20403 ( .A(n21023), .B(n30685), .C(n30636), .Y(n30686) );
  AOI22X1 U20404 ( .A(n25959), .B(n32200), .C(n25791), .D(n23312), .Y(n30692)
         );
  OAI21X1 U20405 ( .A(n25227), .B(n27215), .C(n23145), .Y(n30689) );
  NAND3X1 U20406 ( .A(n24173), .B(n24331), .C(n22817), .Y(n22059) );
  AOI22X1 U20407 ( .A(n26311), .B(n23313), .C(n25988), .D(n32204), .Y(n30700)
         );
  AOI21X1 U20408 ( .A(n29269), .B(n27090), .C(n26282), .Y(n30694) );
  OAI21X1 U20409 ( .A(n23313), .B(n29260), .C(n21928), .Y(n30695) );
  OAI21X1 U20410 ( .A(n32204), .B(n29254), .C(n26326), .Y(n30696) );
  AOI21X1 U20411 ( .A(n26461), .B(n32205), .C(n22158), .Y(n30698) );
  AOI22X1 U20412 ( .A(n21002), .B(n32205), .C(n25555), .D(n23313), .Y(n30705)
         );
  OAI21X1 U20413 ( .A(n30706), .B(n29237), .C(n23002), .Y(n30702) );
  NOR3X1 U20414 ( .A(n30702), .B(n29283), .C(n30701), .Y(n30703) );
  NAND3X1 U20415 ( .A(n24238), .B(n30703), .C(n22736), .Y(n22064) );
  AOI21X1 U20416 ( .A(n29315), .B(n27070), .C(n29280), .Y(n30712) );
  AOI22X1 U20417 ( .A(n25939), .B(n32205), .C(n25790), .D(n23313), .Y(n30711)
         );
  OAI21X1 U20418 ( .A(n25229), .B(n27215), .C(n23147), .Y(n30709) );
  NAND3X1 U20419 ( .A(n24174), .B(n24333), .C(n22818), .Y(n22063) );
  AOI22X1 U20420 ( .A(n26314), .B(n23314), .C(n26037), .D(n32209), .Y(n30720)
         );
  AOI21X1 U20421 ( .A(n29269), .B(n26816), .C(n21056), .Y(n30714) );
  OAI21X1 U20422 ( .A(n23314), .B(n29260), .C(n21929), .Y(n30715) );
  OAI21X1 U20423 ( .A(n32209), .B(n29254), .C(n26328), .Y(n30716) );
  AOI21X1 U20424 ( .A(n26460), .B(n32210), .C(n22162), .Y(n30718) );
  AOI22X1 U20425 ( .A(n29235), .B(n32210), .C(n25535), .D(n23314), .Y(n30725)
         );
  OAI21X1 U20426 ( .A(n30726), .B(n29237), .C(n25185), .Y(n30722) );
  NOR3X1 U20427 ( .A(n30721), .B(n29283), .C(n30722), .Y(n30723) );
  NAND3X1 U20428 ( .A(n30723), .B(n24448), .C(n22737), .Y(n22068) );
  AOI21X1 U20429 ( .A(n29315), .B(n26990), .C(n29277), .Y(n30732) );
  AOI22X1 U20430 ( .A(n25953), .B(n32210), .C(n25799), .D(n23314), .Y(n30731)
         );
  OAI21X1 U20431 ( .A(n25231), .B(n27215), .C(n21040), .Y(n30729) );
  NAND3X1 U20432 ( .A(n24175), .B(n24334), .C(n22819), .Y(n22067) );
  AOI22X1 U20433 ( .A(n26319), .B(n23315), .C(n26036), .D(n32214), .Y(n30739)
         );
  AOI21X1 U20434 ( .A(n29269), .B(n27088), .C(n26303), .Y(n30733) );
  OAI21X1 U20435 ( .A(n23315), .B(n29260), .C(n21930), .Y(n30734) );
  OAI21X1 U20436 ( .A(n32214), .B(n29254), .C(n26330), .Y(n30735) );
  AOI21X1 U20437 ( .A(n26459), .B(n32215), .C(n22166), .Y(n30737) );
  AOI22X1 U20438 ( .A(n20820), .B(n32215), .C(n25534), .D(n23315), .Y(n30744)
         );
  OAI21X1 U20439 ( .A(n30745), .B(n29237), .C(n23003), .Y(n30741) );
  NOR3X1 U20440 ( .A(n30741), .B(n29283), .C(n30740), .Y(n30742) );
  NAND3X1 U20441 ( .A(n30742), .B(n24449), .C(n22738), .Y(n22072) );
  AOI21X1 U20442 ( .A(n29315), .B(n26925), .C(n29277), .Y(n30752) );
  AOI22X1 U20443 ( .A(n25938), .B(n32215), .C(n25789), .D(n23315), .Y(n30751)
         );
  OAI21X1 U20444 ( .A(n25233), .B(n27215), .C(n21047), .Y(n30748) );
  NAND3X1 U20445 ( .A(n24176), .B(n24336), .C(n22820), .Y(n22071) );
  AOI22X1 U20446 ( .A(n26317), .B(n23316), .C(n26004), .D(n32219), .Y(n30760)
         );
  OAI21X1 U20447 ( .A(n23316), .B(n29260), .C(n30754), .Y(n30755) );
  OAI21X1 U20448 ( .A(n32219), .B(n29254), .C(n26328), .Y(n30756) );
  AOI21X1 U20449 ( .A(n26458), .B(n32220), .C(n22169), .Y(n30758) );
  AOI22X1 U20450 ( .A(n20819), .B(n32220), .C(n25537), .D(n23316), .Y(n30765)
         );
  OAI21X1 U20451 ( .A(n30766), .B(n29237), .C(n23004), .Y(n30762) );
  NOR3X1 U20452 ( .A(n29283), .B(n30761), .C(n30762), .Y(n30763) );
  NAND3X1 U20453 ( .A(n24239), .B(n30763), .C(n22739), .Y(n22076) );
  AOI21X1 U20454 ( .A(n29315), .B(n26865), .C(n29277), .Y(n30772) );
  AOI22X1 U20455 ( .A(n25937), .B(n32220), .C(n25791), .D(n23316), .Y(n30771)
         );
  OAI21X1 U20456 ( .A(n25235), .B(n27215), .C(n23151), .Y(n30769) );
  NAND3X1 U20457 ( .A(n24177), .B(n24338), .C(n22821), .Y(n22075) );
  AOI22X1 U20458 ( .A(n26308), .B(n23317), .C(n26039), .D(n32224), .Y(n30779)
         );
  AOI21X1 U20459 ( .A(n29269), .B(n27002), .C(n26299), .Y(n30773) );
  OAI21X1 U20460 ( .A(n23317), .B(n29260), .C(n21931), .Y(n30774) );
  OAI21X1 U20461 ( .A(n32224), .B(n29254), .C(n26327), .Y(n30775) );
  AOI21X1 U20462 ( .A(n26457), .B(n32225), .C(n22170), .Y(n30777) );
  AOI22X1 U20463 ( .A(n20997), .B(n32225), .C(n25549), .D(n23317), .Y(n30784)
         );
  OAI21X1 U20464 ( .A(n30785), .B(n29237), .C(n23005), .Y(n30781) );
  NOR3X1 U20465 ( .A(n30780), .B(n29283), .C(n30781), .Y(n30782) );
  NAND3X1 U20466 ( .A(n24240), .B(n30782), .C(n22740), .Y(n22080) );
  AOI21X1 U20467 ( .A(n29315), .B(n26809), .C(n29277), .Y(n30792) );
  AOI22X1 U20468 ( .A(n25979), .B(n32225), .C(n25786), .D(n23317), .Y(n30791)
         );
  OAI21X1 U20469 ( .A(n25237), .B(n29243), .C(n23153), .Y(n30788) );
  NAND3X1 U20470 ( .A(n24178), .B(n24340), .C(n22822), .Y(n22079) );
  AOI22X1 U20471 ( .A(n26307), .B(n31955), .C(n26011), .D(n32229), .Y(n30800)
         );
  AOI21X1 U20472 ( .A(n29269), .B(n26875), .C(n26280), .Y(n30794) );
  OAI21X1 U20473 ( .A(n31955), .B(n29260), .C(n21932), .Y(n30795) );
  OAI21X1 U20474 ( .A(n32229), .B(n29254), .C(n26323), .Y(n30796) );
  AOI21X1 U20475 ( .A(n26456), .B(n32230), .C(n24034), .Y(n30798) );
  AOI22X1 U20476 ( .A(n29234), .B(n32230), .C(n25553), .D(n31955), .Y(n30805)
         );
  OAI21X1 U20477 ( .A(n30806), .B(n29237), .C(n23006), .Y(n30802) );
  NOR3X1 U20478 ( .A(n30802), .B(n29283), .C(n30801), .Y(n30803) );
  NAND3X1 U20479 ( .A(n24241), .B(n30803), .C(n22741), .Y(n22084) );
  AOI21X1 U20480 ( .A(n29315), .B(n26757), .C(n29277), .Y(n30812) );
  AOI22X1 U20481 ( .A(n25978), .B(n32230), .C(n25796), .D(n31955), .Y(n30811)
         );
  OAI21X1 U20482 ( .A(n25239), .B(n29243), .C(n23117), .Y(n30809) );
  NAND3X1 U20483 ( .A(n24179), .B(n24342), .C(n22823), .Y(n22083) );
  AOI22X1 U20484 ( .A(n26316), .B(n23318), .C(n26038), .D(n32234), .Y(n30819)
         );
  AOI21X1 U20485 ( .A(n29269), .B(n26716), .C(n21078), .Y(n30813) );
  OAI21X1 U20486 ( .A(n23318), .B(n29260), .C(n21933), .Y(n30814) );
  OAI21X1 U20487 ( .A(n32234), .B(n29254), .C(n26331), .Y(n30815) );
  AOI21X1 U20488 ( .A(n26453), .B(n32235), .C(n22174), .Y(n30817) );
  AOI22X1 U20489 ( .A(n20825), .B(n32235), .C(n25555), .D(n23318), .Y(n30824)
         );
  OAI21X1 U20490 ( .A(n30825), .B(n29237), .C(n23007), .Y(n30821) );
  NOR3X1 U20491 ( .A(n29283), .B(n30821), .C(n30820), .Y(n30822) );
  NAND3X1 U20492 ( .A(n24243), .B(n30822), .C(n22742), .Y(n22088) );
  AOI21X1 U20493 ( .A(n29315), .B(n26714), .C(n29278), .Y(n30832) );
  AOI22X1 U20494 ( .A(n25977), .B(n32235), .C(n25787), .D(n23318), .Y(n30831)
         );
  OAI21X1 U20495 ( .A(n25241), .B(n29243), .C(n23155), .Y(n30828) );
  NAND3X1 U20496 ( .A(n24180), .B(n24344), .C(n22824), .Y(n22087) );
  AOI22X1 U20497 ( .A(n26313), .B(n23319), .C(n26042), .D(n32239), .Y(n30840)
         );
  AOI21X1 U20498 ( .A(n29269), .B(n26763), .C(n26297), .Y(n30834) );
  OAI21X1 U20499 ( .A(n23319), .B(n29260), .C(n21934), .Y(n30835) );
  OAI21X1 U20500 ( .A(n32239), .B(n29254), .C(n26334), .Y(n30836) );
  AOI21X1 U20501 ( .A(n26455), .B(n32240), .C(n22177), .Y(n30838) );
  NAND3X1 U20502 ( .A(n24049), .B(n24450), .C(n22796), .Y(n22093) );
  AOI22X1 U20503 ( .A(n29197), .B(n32240), .C(n25568), .D(n23319), .Y(n30845)
         );
  OAI21X1 U20504 ( .A(n30846), .B(n29237), .C(n23008), .Y(n30842) );
  NOR3X1 U20505 ( .A(n30841), .B(n29283), .C(n30842), .Y(n30843) );
  NAND3X1 U20506 ( .A(n21444), .B(n22290), .C(n30843), .Y(n22092) );
  AOI21X1 U20507 ( .A(n29315), .B(n26681), .C(n29277), .Y(n30852) );
  AOI22X1 U20508 ( .A(n25941), .B(n32240), .C(n25788), .D(n23319), .Y(n30851)
         );
  OAI21X1 U20509 ( .A(n25243), .B(n29243), .C(n23191), .Y(n30849) );
  NAND3X1 U20510 ( .A(n24181), .B(n24346), .C(n22825), .Y(n22091) );
  AOI22X1 U20511 ( .A(n26312), .B(n23320), .C(n26009), .D(n32244), .Y(n30859)
         );
  AOI21X1 U20512 ( .A(n29269), .B(n26937), .C(n26284), .Y(n30853) );
  OAI21X1 U20513 ( .A(n23320), .B(n29260), .C(n21935), .Y(n30854) );
  OAI21X1 U20514 ( .A(n32244), .B(n29254), .C(n26324), .Y(n30855) );
  AOI21X1 U20515 ( .A(n26471), .B(n32245), .C(n22178), .Y(n30857) );
  AOI22X1 U20516 ( .A(n20997), .B(n32245), .C(n25545), .D(n23320), .Y(n30864)
         );
  OAI21X1 U20517 ( .A(n30865), .B(n29237), .C(n23192), .Y(n30861) );
  NOR3X1 U20518 ( .A(n30861), .B(n29283), .C(n30860), .Y(n30862) );
  NAND3X1 U20519 ( .A(n24451), .B(n30862), .C(n22294), .Y(n22096) );
  AOI21X1 U20520 ( .A(n29315), .B(n26649), .C(n29280), .Y(n30872) );
  AOI22X1 U20521 ( .A(n25976), .B(n32245), .C(n25787), .D(n23320), .Y(n30871)
         );
  OAI21X1 U20522 ( .A(n25245), .B(n29243), .C(n21038), .Y(n30868) );
  NAND3X1 U20523 ( .A(n24182), .B(n24348), .C(n22826), .Y(n22095) );
  AOI22X1 U20524 ( .A(n26305), .B(n23322), .C(n26041), .D(n32249), .Y(n30880)
         );
  OAI21X1 U20525 ( .A(n23322), .B(n29260), .C(n21989), .Y(n30875) );
  OAI21X1 U20526 ( .A(n32249), .B(n29254), .C(n26330), .Y(n30876) );
  AOI21X1 U20527 ( .A(n26454), .B(n32250), .C(n22182), .Y(n30878) );
  NAND3X1 U20528 ( .A(n22298), .B(n24452), .C(n22797), .Y(n22101) );
  AOI22X1 U20529 ( .A(n29197), .B(n32250), .C(n25554), .D(n23322), .Y(n30885)
         );
  OAI21X1 U20530 ( .A(n30886), .B(n29237), .C(n23009), .Y(n30882) );
  NOR3X1 U20531 ( .A(n30882), .B(n29283), .C(n30881), .Y(n30883) );
  NAND3X1 U20532 ( .A(n22302), .B(n24453), .C(n30883), .Y(n22100) );
  AOI21X1 U20533 ( .A(n29315), .B(n26623), .C(n29278), .Y(n30893) );
  AOI22X1 U20534 ( .A(n25975), .B(n32250), .C(n25786), .D(n23322), .Y(n30892)
         );
  OAI21X1 U20535 ( .A(n25247), .B(n27215), .C(n23077), .Y(n30889) );
  NAND3X1 U20536 ( .A(n24183), .B(n24350), .C(n22827), .Y(n22099) );
  AOI22X1 U20537 ( .A(n26310), .B(n23323), .C(n25986), .D(n32254), .Y(n30900)
         );
  OAI21X1 U20538 ( .A(n23323), .B(n29261), .C(n30894), .Y(n30895) );
  OAI21X1 U20539 ( .A(n32254), .B(n29255), .C(n26324), .Y(n30896) );
  AOI21X1 U20540 ( .A(n26469), .B(n32255), .C(n24035), .Y(n30898) );
  NAND3X1 U20541 ( .A(n22653), .B(n24454), .C(n24051), .Y(n22105) );
  AOI22X1 U20542 ( .A(n29197), .B(n32255), .C(n25540), .D(n23323), .Y(n30905)
         );
  OAI21X1 U20543 ( .A(n30906), .B(n29238), .C(n23010), .Y(n30902) );
  NOR3X1 U20544 ( .A(n30902), .B(n29283), .C(n30901), .Y(n30903) );
  NAND3X1 U20545 ( .A(n22306), .B(n24455), .C(n30903), .Y(n22104) );
  AOI21X1 U20546 ( .A(n29316), .B(n27165), .C(n29280), .Y(n30913) );
  AOI22X1 U20547 ( .A(n25947), .B(n32255), .C(n25790), .D(n23323), .Y(n30912)
         );
  OAI21X1 U20548 ( .A(n25249), .B(n29243), .C(n23134), .Y(n30909) );
  NAND3X1 U20549 ( .A(n24184), .B(n24352), .C(n22828), .Y(n22103) );
  AOI22X1 U20550 ( .A(n26316), .B(n23324), .C(n25984), .D(n32259), .Y(n30921)
         );
  AOI21X1 U20551 ( .A(n29268), .B(n26818), .C(n26298), .Y(n30915) );
  OAI21X1 U20552 ( .A(n23324), .B(n29261), .C(n21936), .Y(n30916) );
  OAI21X1 U20553 ( .A(n32259), .B(n29255), .C(n26324), .Y(n30917) );
  AOI21X1 U20554 ( .A(n26466), .B(n32260), .C(n24036), .Y(n30919) );
  AOI22X1 U20555 ( .A(n29235), .B(n32260), .C(n25553), .D(n23324), .Y(n30926)
         );
  OAI21X1 U20556 ( .A(n30927), .B(n29238), .C(n23011), .Y(n30923) );
  NOR3X1 U20557 ( .A(n30923), .B(n29284), .C(n30922), .Y(n30924) );
  NAND3X1 U20558 ( .A(n24456), .B(n22307), .C(n30924), .Y(n22108) );
  AOI21X1 U20559 ( .A(n29315), .B(n27069), .C(n29278), .Y(n30933) );
  AOI22X1 U20560 ( .A(n25955), .B(n32260), .C(n25797), .D(n23324), .Y(n30932)
         );
  OAI21X1 U20561 ( .A(n25251), .B(n25856), .C(n21046), .Y(n30930) );
  NAND3X1 U20562 ( .A(n24185), .B(n24354), .C(n22829), .Y(n22107) );
  AOI22X1 U20563 ( .A(n26320), .B(n32266), .C(n25985), .D(n32264), .Y(n30940)
         );
  AOI21X1 U20564 ( .A(n29268), .B(n27094), .C(n21078), .Y(n30934) );
  OAI21X1 U20565 ( .A(n32264), .B(n29255), .C(n26324), .Y(n30936) );
  AOI21X1 U20566 ( .A(n26460), .B(n32265), .C(n22190), .Y(n30938) );
  AOI22X1 U20567 ( .A(n29235), .B(n32265), .C(n25542), .D(n32266), .Y(n30945)
         );
  OAI21X1 U20568 ( .A(n30946), .B(n29238), .C(n23012), .Y(n30942) );
  NOR3X1 U20569 ( .A(n30942), .B(n29284), .C(n30941), .Y(n30943) );
  NAND3X1 U20570 ( .A(n22310), .B(n24457), .C(n30943), .Y(n22112) );
  AOI21X1 U20571 ( .A(n29316), .B(n26924), .C(n29278), .Y(n30953) );
  AOI22X1 U20572 ( .A(n25954), .B(n32265), .C(n25797), .D(n32266), .Y(n30952)
         );
  OAI21X1 U20573 ( .A(n25253), .B(n29244), .C(n23193), .Y(n30949) );
  NAND3X1 U20574 ( .A(n24186), .B(n24356), .C(n22830), .Y(n22111) );
  AOI22X1 U20575 ( .A(n26316), .B(n23325), .C(n26007), .D(n32270), .Y(n30961)
         );
  AOI21X1 U20576 ( .A(n29268), .B(n27092), .C(n20839), .Y(n30955) );
  OAI21X1 U20577 ( .A(n23325), .B(n29261), .C(n21937), .Y(n30956) );
  OAI21X1 U20578 ( .A(n32270), .B(n29255), .C(n26324), .Y(n30957) );
  AOI21X1 U20579 ( .A(n26470), .B(n32271), .C(n24037), .Y(n30959) );
  NAND3X1 U20580 ( .A(n24053), .B(n24458), .C(n22798), .Y(n22117) );
  AOI22X1 U20581 ( .A(n29235), .B(n32271), .C(n25554), .D(n23325), .Y(n30966)
         );
  OAI21X1 U20582 ( .A(n30967), .B(n29238), .C(n23013), .Y(n30963) );
  NOR3X1 U20583 ( .A(n30963), .B(n29284), .C(n30962), .Y(n30964) );
  NAND3X1 U20584 ( .A(n22311), .B(n24459), .C(n30964), .Y(n22116) );
  AOI21X1 U20585 ( .A(n29316), .B(n26989), .C(n29278), .Y(n30974) );
  AOI22X1 U20586 ( .A(n25941), .B(n32271), .C(n25789), .D(n23325), .Y(n30973)
         );
  OAI21X1 U20587 ( .A(n25255), .B(n25856), .C(n23121), .Y(n30970) );
  NAND3X1 U20588 ( .A(n24187), .B(n24358), .C(n22831), .Y(n22115) );
  AOI22X1 U20589 ( .A(n26315), .B(n23328), .C(n25987), .D(n32275), .Y(n30982)
         );
  AOI21X1 U20590 ( .A(n29268), .B(n25358), .C(n20839), .Y(n30976) );
  OAI21X1 U20591 ( .A(n23328), .B(n29261), .C(n21938), .Y(n30977) );
  OAI21X1 U20592 ( .A(n32275), .B(n29255), .C(n26335), .Y(n30978) );
  AOI21X1 U20593 ( .A(n26468), .B(n23327), .C(n22198), .Y(n30980) );
  NAND3X1 U20594 ( .A(n22312), .B(n24460), .C(n24850), .Y(n22121) );
  AOI22X1 U20595 ( .A(n29235), .B(n23327), .C(n25550), .D(n23328), .Y(n30986)
         );
  OAI21X1 U20596 ( .A(n30987), .B(n29238), .C(n23014), .Y(n30983) );
  NOR3X1 U20597 ( .A(n30983), .B(n29284), .C(n30989), .Y(n30984) );
  NAND3X1 U20598 ( .A(n22313), .B(n24461), .C(n30984), .Y(n22120) );
  AOI21X1 U20599 ( .A(n29316), .B(n26864), .C(n29278), .Y(n30994) );
  AOI22X1 U20600 ( .A(n25974), .B(n23327), .C(n25788), .D(n23328), .Y(n30993)
         );
  OAI21X1 U20601 ( .A(n25257), .B(n25757), .C(n25652), .Y(n30990) );
  NAND3X1 U20602 ( .A(n24188), .B(n24360), .C(n22832), .Y(n22119) );
  AOI22X1 U20603 ( .A(n26478), .B(n32279), .C(n26310), .D(n23330), .Y(n31000)
         );
  OAI21X1 U20604 ( .A(n23329), .B(n29255), .C(n26326), .Y(n30995) );
  OAI21X1 U20605 ( .A(n23330), .B(n29261), .C(n30996), .Y(n30997) );
  NOR3X1 U20606 ( .A(n27230), .B(n31851), .C(n31006), .Y(n30998) );
  NAND3X1 U20607 ( .A(n30998), .B(n24462), .C(n22314), .Y(n22125) );
  AOI22X1 U20608 ( .A(n25545), .B(n23330), .C(n25892), .D(n23329), .Y(n31005)
         );
  NOR3X1 U20609 ( .A(n31006), .B(n29277), .C(n31002), .Y(n31003) );
  NAND3X1 U20610 ( .A(n24055), .B(n24463), .C(n31003), .Y(n22124) );
  AOI21X1 U20611 ( .A(n25950), .B(n32279), .C(n29287), .Y(n31010) );
  AOI22X1 U20612 ( .A(n25815), .B(n23330), .C(n25854), .D(n23329), .Y(n31009)
         );
  OAI21X1 U20613 ( .A(n31001), .B(n27146), .C(n23015), .Y(n31007) );
  NAND3X1 U20614 ( .A(n24189), .B(n24362), .C(n22833), .Y(n22123) );
  AOI22X1 U20615 ( .A(n26315), .B(n23333), .C(n26006), .D(n32283), .Y(n31018)
         );
  AOI21X1 U20616 ( .A(n29268), .B(n25359), .C(n26284), .Y(n31012) );
  OAI21X1 U20617 ( .A(n23333), .B(n29261), .C(n21939), .Y(n31013) );
  OAI21X1 U20618 ( .A(n32283), .B(n29255), .C(n26324), .Y(n31014) );
  AOI21X1 U20619 ( .A(n26462), .B(n23332), .C(n22206), .Y(n31016) );
  AOI22X1 U20620 ( .A(n29234), .B(n23332), .C(n25551), .D(n23333), .Y(n31023)
         );
  OAI21X1 U20621 ( .A(n31024), .B(n29238), .C(n23195), .Y(n31020) );
  NOR3X1 U20622 ( .A(n29284), .B(n31020), .C(n31019), .Y(n31021) );
  NAND3X1 U20623 ( .A(n22315), .B(n24464), .C(n31021), .Y(n22128) );
  AOI21X1 U20624 ( .A(n29316), .B(n26808), .C(n29278), .Y(n31031) );
  AOI22X1 U20625 ( .A(n25970), .B(n23332), .C(n25796), .D(n23333), .Y(n31030)
         );
  OAI21X1 U20626 ( .A(n25259), .B(n25758), .C(n23158), .Y(n31027) );
  NAND3X1 U20627 ( .A(n24190), .B(n24364), .C(n22834), .Y(n22127) );
  AOI22X1 U20628 ( .A(n21004), .B(n32287), .C(n26318), .D(n23335), .Y(n31037)
         );
  OAI21X1 U20629 ( .A(n23334), .B(n29255), .C(n26334), .Y(n31032) );
  AOI21X1 U20630 ( .A(n29268), .B(n26759), .C(n26290), .Y(n31033) );
  OAI21X1 U20631 ( .A(n23335), .B(n29261), .C(n21940), .Y(n31034) );
  NOR3X1 U20632 ( .A(n27231), .B(n31897), .C(n31039), .Y(n31035) );
  NAND3X1 U20633 ( .A(n24465), .B(n31035), .C(n22316), .Y(n22133) );
  AOI22X1 U20634 ( .A(n25547), .B(n23335), .C(n25893), .D(n23334), .Y(n31043)
         );
  NOR3X1 U20635 ( .A(n31040), .B(n29280), .C(n31039), .Y(n31041) );
  NAND3X1 U20636 ( .A(n24057), .B(n24466), .C(n31041), .Y(n22132) );
  AOI21X1 U20637 ( .A(n25951), .B(n32287), .C(n29287), .Y(n31048) );
  AOI22X1 U20638 ( .A(n25816), .B(n23335), .C(n25854), .D(n23334), .Y(n31047)
         );
  OAI21X1 U20639 ( .A(n31038), .B(n27146), .C(n23016), .Y(n31045) );
  NAND3X1 U20640 ( .A(n24191), .B(n24366), .C(n22835), .Y(n22131) );
  AOI22X1 U20641 ( .A(n26305), .B(n23337), .C(n26005), .D(n32291), .Y(n31056)
         );
  OAI21X1 U20642 ( .A(n23337), .B(n29261), .C(n31050), .Y(n31051) );
  OAI21X1 U20643 ( .A(n32291), .B(n29255), .C(n26324), .Y(n31052) );
  AOI21X1 U20644 ( .A(n26477), .B(n23336), .C(n22214), .Y(n31054) );
  NAND3X1 U20645 ( .A(n23607), .B(n24467), .C(n22799), .Y(n22137) );
  AOI22X1 U20646 ( .A(n20827), .B(n23336), .C(n25552), .D(n23337), .Y(n31061)
         );
  OAI21X1 U20647 ( .A(n31062), .B(n29238), .C(n23018), .Y(n31058) );
  NOR3X1 U20648 ( .A(n31058), .B(n29284), .C(n31057), .Y(n31059) );
  NAND3X1 U20649 ( .A(n22317), .B(n24468), .C(n31059), .Y(n22136) );
  AOI21X1 U20650 ( .A(n29316), .B(n26756), .C(n29278), .Y(n31069) );
  AOI22X1 U20651 ( .A(n25970), .B(n23336), .C(n25795), .D(n23337), .Y(n31068)
         );
  OAI21X1 U20652 ( .A(n25260), .B(n25757), .C(n23160), .Y(n31065) );
  NAND3X1 U20653 ( .A(n24192), .B(n24368), .C(n22836), .Y(n22135) );
  AOI22X1 U20654 ( .A(n26448), .B(n32295), .C(n26313), .D(n23339), .Y(n31075)
         );
  OAI21X1 U20655 ( .A(n23338), .B(n29255), .C(n26335), .Y(n31070) );
  AOI21X1 U20656 ( .A(n29268), .B(n27111), .C(n26282), .Y(n31071) );
  OAI21X1 U20657 ( .A(n23339), .B(n29261), .C(n21941), .Y(n31072) );
  NOR3X1 U20658 ( .A(n31085), .B(n31897), .C(n31078), .Y(n31073) );
  NAND3X1 U20659 ( .A(n31073), .B(n24469), .C(n22318), .Y(n22141) );
  AOI22X1 U20660 ( .A(n25543), .B(n23339), .C(n25894), .D(n23338), .Y(n31082)
         );
  OAI21X1 U20661 ( .A(n27110), .B(n29208), .C(n26972), .Y(n31079) );
  NOR3X1 U20662 ( .A(n29277), .B(n31079), .C(n31078), .Y(n31080) );
  NAND3X1 U20663 ( .A(n22319), .B(n24470), .C(n31080), .Y(n22140) );
  AOI21X1 U20664 ( .A(n25948), .B(n32295), .C(n29287), .Y(n31088) );
  AOI22X1 U20665 ( .A(n25815), .B(n23339), .C(n25854), .D(n23338), .Y(n31087)
         );
  OAI21X1 U20666 ( .A(n31076), .B(n27146), .C(n23019), .Y(n31084) );
  NAND3X1 U20667 ( .A(n24193), .B(n24370), .C(n22837), .Y(n22139) );
  AOI22X1 U20668 ( .A(n26314), .B(n23341), .C(n26011), .D(n32299), .Y(n31096)
         );
  AOI21X1 U20669 ( .A(n29268), .B(n25361), .C(n26303), .Y(n31090) );
  OAI21X1 U20670 ( .A(n23341), .B(n29261), .C(n21942), .Y(n31091) );
  OAI21X1 U20671 ( .A(n32299), .B(n29255), .C(n26324), .Y(n31092) );
  AOI21X1 U20672 ( .A(n26479), .B(n23340), .C(n22222), .Y(n31094) );
  AOI22X1 U20673 ( .A(n21003), .B(n23340), .C(n25565), .D(n23341), .Y(n31101)
         );
  OAI21X1 U20674 ( .A(n31102), .B(n29238), .C(n23196), .Y(n31098) );
  NOR3X1 U20675 ( .A(n29284), .B(n31098), .C(n31097), .Y(n31099) );
  NAND3X1 U20676 ( .A(n31099), .B(n23459), .C(n22320), .Y(n22144) );
  AOI21X1 U20677 ( .A(n29316), .B(n26713), .C(n29278), .Y(n31109) );
  AOI22X1 U20678 ( .A(n25969), .B(n23340), .C(n25795), .D(n23341), .Y(n31108)
         );
  OAI21X1 U20679 ( .A(n25262), .B(n29244), .C(n23162), .Y(n31105) );
  NAND3X1 U20680 ( .A(n24194), .B(n24372), .C(n22838), .Y(n22143) );
  AOI22X1 U20681 ( .A(n26473), .B(n32303), .C(n26307), .D(n23343), .Y(n31115)
         );
  OAI21X1 U20682 ( .A(n23342), .B(n29255), .C(n26324), .Y(n31110) );
  AOI21X1 U20683 ( .A(n29268), .B(n27014), .C(n26283), .Y(n31111) );
  OAI21X1 U20684 ( .A(n23343), .B(n29261), .C(n21943), .Y(n31112) );
  NOR3X1 U20685 ( .A(n31125), .B(n31897), .C(n31118), .Y(n31113) );
  NAND3X1 U20686 ( .A(n22321), .B(n24471), .C(n31113), .Y(n22149) );
  AOI22X1 U20687 ( .A(n25546), .B(n23343), .C(n25891), .D(n23342), .Y(n31122)
         );
  OAI21X1 U20688 ( .A(n27013), .B(n29236), .C(n23020), .Y(n31119) );
  NOR3X1 U20689 ( .A(n29277), .B(n31119), .C(n31118), .Y(n31120) );
  NAND3X1 U20690 ( .A(n22322), .B(n24472), .C(n31120), .Y(n22148) );
  AOI21X1 U20691 ( .A(n25945), .B(n32303), .C(n29287), .Y(n31128) );
  AOI22X1 U20692 ( .A(n25816), .B(n23343), .C(n25854), .D(n23342), .Y(n31127)
         );
  OAI21X1 U20693 ( .A(n31116), .B(n27146), .C(n23021), .Y(n31124) );
  NAND3X1 U20694 ( .A(n24195), .B(n24374), .C(n22839), .Y(n22147) );
  AOI22X1 U20695 ( .A(n26320), .B(n23345), .C(n26008), .D(n32307), .Y(n31136)
         );
  AOI21X1 U20696 ( .A(n29268), .B(n25362), .C(n20840), .Y(n31130) );
  OAI21X1 U20697 ( .A(n23345), .B(n29261), .C(n21944), .Y(n31131) );
  OAI21X1 U20698 ( .A(n32307), .B(n29256), .C(n26324), .Y(n31132) );
  AOI21X1 U20699 ( .A(n26467), .B(n23344), .C(n24038), .Y(n31134) );
  NAND3X1 U20700 ( .A(n24059), .B(n24473), .C(n22800), .Y(n22153) );
  AOI22X1 U20701 ( .A(n20824), .B(n23344), .C(n25552), .D(n23345), .Y(n31141)
         );
  OAI21X1 U20702 ( .A(n31142), .B(n29238), .C(n23023), .Y(n31138) );
  NOR3X1 U20703 ( .A(n31138), .B(n29284), .C(n31137), .Y(n31139) );
  NAND3X1 U20704 ( .A(n22375), .B(n24474), .C(n31139), .Y(n22152) );
  AOI21X1 U20705 ( .A(n29316), .B(n26680), .C(n29278), .Y(n31149) );
  AOI22X1 U20706 ( .A(n25968), .B(n23344), .C(n25794), .D(n23345), .Y(n31148)
         );
  OAI21X1 U20707 ( .A(n25264), .B(n29244), .C(n23122), .Y(n31145) );
  NAND3X1 U20708 ( .A(n24196), .B(n24376), .C(n22840), .Y(n22151) );
  AOI22X1 U20709 ( .A(n26468), .B(n32311), .C(n26319), .D(n23456), .Y(n31155)
         );
  OAI21X1 U20710 ( .A(n23346), .B(n29256), .C(n26327), .Y(n31150) );
  NOR3X1 U20711 ( .A(n27228), .B(n31897), .C(n31157), .Y(n31153) );
  NAND3X1 U20712 ( .A(n24475), .B(n22420), .C(n31153), .Y(n22157) );
  AOI22X1 U20713 ( .A(n25547), .B(n23456), .C(n25898), .D(n23346), .Y(n31161)
         );
  NOR3X1 U20714 ( .A(n29277), .B(n31158), .C(n31157), .Y(n31159) );
  NAND3X1 U20715 ( .A(n24061), .B(n24476), .C(n31159), .Y(n22156) );
  AOI21X1 U20716 ( .A(n25948), .B(n32311), .C(n29287), .Y(n31166) );
  AOI22X1 U20717 ( .A(n25800), .B(n23456), .C(n25854), .D(n23346), .Y(n31165)
         );
  OAI21X1 U20718 ( .A(n31156), .B(n27146), .C(n20841), .Y(n31163) );
  NAND3X1 U20719 ( .A(n24197), .B(n24378), .C(n22841), .Y(n22155) );
  AOI22X1 U20720 ( .A(n26317), .B(n23348), .C(n26010), .D(n32315), .Y(n31174)
         );
  OAI21X1 U20721 ( .A(n23348), .B(n29261), .C(n21990), .Y(n31169) );
  OAI21X1 U20722 ( .A(n32315), .B(n29256), .C(n26324), .Y(n31170) );
  AOI21X1 U20723 ( .A(n26476), .B(n23347), .C(n22229), .Y(n31172) );
  NAND3X1 U20724 ( .A(n24063), .B(n23460), .C(n22801), .Y(n22161) );
  AOI22X1 U20725 ( .A(n21001), .B(n23347), .C(n25551), .D(n23348), .Y(n31178)
         );
  OAI21X1 U20726 ( .A(n31179), .B(n29238), .C(n23025), .Y(n31175) );
  NOR3X1 U20727 ( .A(n31175), .B(n29284), .C(n25596), .Y(n31176) );
  NAND3X1 U20728 ( .A(n22421), .B(n24477), .C(n31176), .Y(n22160) );
  AOI21X1 U20729 ( .A(n29316), .B(n26648), .C(n29278), .Y(n31186) );
  AOI22X1 U20730 ( .A(n25950), .B(n23347), .C(n25794), .D(n23348), .Y(n31185)
         );
  OAI21X1 U20731 ( .A(n25266), .B(n29246), .C(n23089), .Y(n31182) );
  NAND3X1 U20732 ( .A(n24198), .B(n24380), .C(n22842), .Y(n22159) );
  AOI22X1 U20733 ( .A(n26469), .B(n32319), .C(n26320), .D(n23350), .Y(n31192)
         );
  OAI21X1 U20734 ( .A(n23349), .B(n29256), .C(n26329), .Y(n31187) );
  AOI21X1 U20735 ( .A(n29267), .B(n27108), .C(n26302), .Y(n31188) );
  OAI21X1 U20736 ( .A(n23350), .B(n29261), .C(n21945), .Y(n31189) );
  NOR3X1 U20737 ( .A(n31202), .B(n31851), .C(n31195), .Y(n31190) );
  NAND3X1 U20738 ( .A(n31190), .B(n24478), .C(n22422), .Y(n22165) );
  AOI22X1 U20739 ( .A(n25546), .B(n23350), .C(n25899), .D(n23349), .Y(n31199)
         );
  OAI21X1 U20740 ( .A(n27107), .B(n29208), .C(n26973), .Y(n31196) );
  NOR3X1 U20741 ( .A(n29277), .B(n31196), .C(n31195), .Y(n31197) );
  NAND3X1 U20742 ( .A(n22423), .B(n24479), .C(n31197), .Y(n22164) );
  AOI21X1 U20743 ( .A(n25946), .B(n32319), .C(n29287), .Y(n31205) );
  AOI22X1 U20744 ( .A(n25801), .B(n23350), .C(n25854), .D(n23349), .Y(n31204)
         );
  OAI21X1 U20745 ( .A(n31193), .B(n27146), .C(n23026), .Y(n31201) );
  NAND3X1 U20746 ( .A(n24199), .B(n24382), .C(n22843), .Y(n22163) );
  AOI22X1 U20747 ( .A(n26313), .B(n23352), .C(n26012), .D(n32323), .Y(n31213)
         );
  AOI21X1 U20748 ( .A(n29268), .B(n25363), .C(n26287), .Y(n31207) );
  OAI21X1 U20749 ( .A(n23352), .B(n29261), .C(n21946), .Y(n31208) );
  OAI21X1 U20750 ( .A(n32323), .B(n29256), .C(n26327), .Y(n31209) );
  AOI21X1 U20751 ( .A(n26466), .B(n23351), .C(n22230), .Y(n31211) );
  AOI22X1 U20752 ( .A(n20829), .B(n23351), .C(n25536), .D(n23352), .Y(n31218)
         );
  OAI21X1 U20753 ( .A(n31219), .B(n29238), .C(n23028), .Y(n31215) );
  NOR3X1 U20754 ( .A(n31215), .B(n29284), .C(n31214), .Y(n31216) );
  NAND3X1 U20755 ( .A(n31216), .B(n21447), .C(n22743), .Y(n22168) );
  AOI21X1 U20756 ( .A(n29316), .B(n26622), .C(n29278), .Y(n31226) );
  AOI22X1 U20757 ( .A(n25967), .B(n23351), .C(n25823), .D(n23352), .Y(n31225)
         );
  OAI21X1 U20758 ( .A(n25268), .B(n25757), .C(n23164), .Y(n31222) );
  NAND3X1 U20759 ( .A(n24200), .B(n24384), .C(n22844), .Y(n22167) );
  AOI22X1 U20760 ( .A(n26470), .B(n32327), .C(n26307), .D(n23354), .Y(n31232)
         );
  OAI21X1 U20761 ( .A(n23353), .B(n29256), .C(n26324), .Y(n31227) );
  AOI21X1 U20762 ( .A(n29269), .B(n27011), .C(n26299), .Y(n31228) );
  OAI21X1 U20763 ( .A(n23354), .B(n29261), .C(n21947), .Y(n31229) );
  NOR3X1 U20764 ( .A(n31242), .B(n31897), .C(n31235), .Y(n31230) );
  NAND3X1 U20765 ( .A(n31230), .B(n24480), .C(n22424), .Y(n22173) );
  AOI22X1 U20766 ( .A(n25544), .B(n23354), .C(n25900), .D(n23353), .Y(n31239)
         );
  OAI21X1 U20767 ( .A(n27010), .B(n29236), .C(n23029), .Y(n31236) );
  NOR3X1 U20768 ( .A(n29277), .B(n31236), .C(n31235), .Y(n31237) );
  NAND3X1 U20769 ( .A(n24065), .B(n24481), .C(n31237), .Y(n22172) );
  AOI21X1 U20770 ( .A(n25947), .B(n32327), .C(n29287), .Y(n31245) );
  AOI22X1 U20771 ( .A(n25802), .B(n23354), .C(n25854), .D(n23353), .Y(n31244)
         );
  OAI21X1 U20772 ( .A(n31233), .B(n27146), .C(n23031), .Y(n31241) );
  NAND3X1 U20773 ( .A(n24201), .B(n24385), .C(n22845), .Y(n22171) );
  AOI22X1 U20774 ( .A(n26312), .B(n23356), .C(n26013), .D(n32331), .Y(n31253)
         );
  AOI21X1 U20775 ( .A(n29266), .B(n25364), .C(n26291), .Y(n31247) );
  OAI21X1 U20776 ( .A(n23356), .B(n29261), .C(n21948), .Y(n31248) );
  OAI21X1 U20777 ( .A(n32331), .B(n29256), .C(n26327), .Y(n31249) );
  AOI21X1 U20778 ( .A(n26479), .B(n23355), .C(n22237), .Y(n31251) );
  AOI22X1 U20779 ( .A(n29232), .B(n23355), .C(n25535), .D(n23356), .Y(n31258)
         );
  OAI21X1 U20780 ( .A(n31259), .B(n29238), .C(n23032), .Y(n31255) );
  NOR3X1 U20781 ( .A(n31255), .B(n29284), .C(n31254), .Y(n31256) );
  NAND3X1 U20782 ( .A(n31256), .B(n21450), .C(n22744), .Y(n22176) );
  AOI21X1 U20783 ( .A(n29316), .B(n26597), .C(n29278), .Y(n31266) );
  AOI22X1 U20784 ( .A(n25966), .B(n23355), .C(n25824), .D(n23356), .Y(n31265)
         );
  OAI21X1 U20785 ( .A(n25270), .B(n25856), .C(n23166), .Y(n31262) );
  NAND3X1 U20786 ( .A(n24202), .B(n24387), .C(n22846), .Y(n22175) );
  AOI22X1 U20787 ( .A(n26449), .B(n32335), .C(n26312), .D(n23357), .Y(n31272)
         );
  OAI21X1 U20788 ( .A(n26275), .B(n29256), .C(n26324), .Y(n31267) );
  AOI21X1 U20789 ( .A(n29267), .B(n26946), .C(n20843), .Y(n31268) );
  OAI21X1 U20790 ( .A(n23357), .B(n29261), .C(n21949), .Y(n31269) );
  NOR3X1 U20791 ( .A(n31274), .B(n31897), .C(n31275), .Y(n31270) );
  NAND3X1 U20792 ( .A(n22434), .B(n24482), .C(n31270), .Y(n22181) );
  AOI22X1 U20793 ( .A(n25540), .B(n23357), .C(n25901), .D(n26275), .Y(n31279)
         );
  OAI21X1 U20794 ( .A(n26945), .B(n29208), .C(n23033), .Y(n31276) );
  NOR3X1 U20795 ( .A(n29277), .B(n31276), .C(n31275), .Y(n31277) );
  NAND3X1 U20796 ( .A(n24067), .B(n24483), .C(n31277), .Y(n22180) );
  AOI21X1 U20797 ( .A(n25943), .B(n32335), .C(n29287), .Y(n31284) );
  AOI22X1 U20798 ( .A(n25803), .B(n23357), .C(n25854), .D(n21169), .Y(n31283)
         );
  OAI21X1 U20799 ( .A(n31273), .B(n27146), .C(n20844), .Y(n31281) );
  NAND3X1 U20800 ( .A(n24203), .B(n24388), .C(n22847), .Y(n22179) );
  AOI22X1 U20801 ( .A(n26311), .B(n23359), .C(n26014), .D(n32339), .Y(n31291)
         );
  AOI21X1 U20802 ( .A(n29269), .B(n25365), .C(n20840), .Y(n31285) );
  OAI21X1 U20803 ( .A(n23359), .B(n29261), .C(n21950), .Y(n31286) );
  OAI21X1 U20804 ( .A(n32339), .B(n29256), .C(n26326), .Y(n31287) );
  AOI21X1 U20805 ( .A(n26478), .B(n23358), .C(n24039), .Y(n31289) );
  NAND3X1 U20806 ( .A(n24069), .B(n24484), .C(n22802), .Y(n22185) );
  AOI22X1 U20807 ( .A(n29235), .B(n23358), .C(n25567), .D(n23359), .Y(n31295)
         );
  OAI21X1 U20808 ( .A(n31296), .B(n29239), .C(n25178), .Y(n31292) );
  NOR3X1 U20809 ( .A(n20833), .B(n29284), .C(n31292), .Y(n31293) );
  NAND3X1 U20810 ( .A(n22437), .B(n21453), .C(n31293), .Y(n22184) );
  AOI21X1 U20811 ( .A(n29316), .B(n27164), .C(n29278), .Y(n31302) );
  AOI22X1 U20812 ( .A(n25965), .B(n23358), .C(n25800), .D(n23359), .Y(n31301)
         );
  OAI21X1 U20813 ( .A(n25272), .B(n29245), .C(n23082), .Y(n31299) );
  NAND3X1 U20814 ( .A(n24204), .B(n24390), .C(n22848), .Y(n22183) );
  AOI22X1 U20815 ( .A(n26310), .B(n23361), .C(n26022), .D(n32343), .Y(n31310)
         );
  OAI21X1 U20816 ( .A(n23361), .B(n29261), .C(n31304), .Y(n31305) );
  OAI21X1 U20817 ( .A(n32343), .B(n29256), .C(n26335), .Y(n31306) );
  AOI21X1 U20818 ( .A(n26478), .B(n23360), .C(n24040), .Y(n31308) );
  NAND3X1 U20819 ( .A(n24070), .B(n24485), .C(n22803), .Y(n22189) );
  AOI22X1 U20820 ( .A(n29197), .B(n23360), .C(n25538), .D(n23361), .Y(n31314)
         );
  OAI21X1 U20821 ( .A(n31315), .B(n29239), .C(n23035), .Y(n31311) );
  NOR3X1 U20822 ( .A(n25515), .B(n29285), .C(n31311), .Y(n31312) );
  NAND3X1 U20823 ( .A(n21456), .B(n22440), .C(n31312), .Y(n22188) );
  AOI21X1 U20824 ( .A(n29317), .B(n27068), .C(n29278), .Y(n31320) );
  AOI22X1 U20825 ( .A(n25951), .B(n23360), .C(n25793), .D(n23361), .Y(n31319)
         );
  OAI21X1 U20826 ( .A(n25274), .B(n25857), .C(n23084), .Y(n31317) );
  NAND3X1 U20827 ( .A(n24205), .B(n24392), .C(n22849), .Y(n22187) );
  AOI22X1 U20828 ( .A(n26314), .B(n23363), .C(n26023), .D(n32347), .Y(n31327)
         );
  AOI21X1 U20829 ( .A(n29269), .B(n25367), .C(n26293), .Y(n31321) );
  OAI21X1 U20830 ( .A(n23363), .B(n29261), .C(n21951), .Y(n31322) );
  OAI21X1 U20831 ( .A(n32347), .B(n29256), .C(n26335), .Y(n31323) );
  AOI21X1 U20832 ( .A(n26474), .B(n23362), .C(n22238), .Y(n31325) );
  NAND3X1 U20833 ( .A(n24071), .B(n24486), .C(n22804), .Y(n22193) );
  AOI22X1 U20834 ( .A(n29235), .B(n23362), .C(n25568), .D(n23363), .Y(n31332)
         );
  OAI21X1 U20835 ( .A(n31333), .B(n29239), .C(n23036), .Y(n31329) );
  NOR3X1 U20836 ( .A(n31328), .B(n29285), .C(n31329), .Y(n31330) );
  NAND3X1 U20837 ( .A(n22443), .B(n21459), .C(n31330), .Y(n22192) );
  AOI21X1 U20838 ( .A(n29317), .B(n26988), .C(n29279), .Y(n31339) );
  AOI22X1 U20839 ( .A(n25964), .B(n23362), .C(n25785), .D(n23363), .Y(n31338)
         );
  OAI21X1 U20840 ( .A(n25276), .B(n29244), .C(n23198), .Y(n31336) );
  NAND3X1 U20841 ( .A(n24206), .B(n24394), .C(n22850), .Y(n22191) );
  AOI22X1 U20842 ( .A(n26310), .B(n23366), .C(n26024), .D(n32351), .Y(n31347)
         );
  OAI21X1 U20843 ( .A(n23366), .B(n29261), .C(n31341), .Y(n31342) );
  OAI21X1 U20844 ( .A(n32351), .B(n29256), .C(n26329), .Y(n31343) );
  AOI21X1 U20845 ( .A(n26477), .B(n23365), .C(n24041), .Y(n31345) );
  NAND3X1 U20846 ( .A(n24072), .B(n24487), .C(n22805), .Y(n22197) );
  AOI22X1 U20847 ( .A(n29235), .B(n23365), .C(n25565), .D(n23366), .Y(n31352)
         );
  OAI21X1 U20848 ( .A(n31353), .B(n29239), .C(n23037), .Y(n31349) );
  NOR3X1 U20849 ( .A(n31349), .B(n29285), .C(n31348), .Y(n31350) );
  NAND3X1 U20850 ( .A(n22446), .B(n21462), .C(n31350), .Y(n22196) );
  AOI21X1 U20851 ( .A(n29317), .B(n26923), .C(n29279), .Y(n31360) );
  AOI22X1 U20852 ( .A(n25963), .B(n23365), .C(n25788), .D(n23366), .Y(n31359)
         );
  OAI21X1 U20853 ( .A(n25278), .B(n25856), .C(n23124), .Y(n31356) );
  NAND3X1 U20854 ( .A(n24207), .B(n24396), .C(n22851), .Y(n22195) );
  AOI22X1 U20855 ( .A(n26322), .B(n23368), .C(n26025), .D(n32355), .Y(n31367)
         );
  AOI21X1 U20856 ( .A(n29267), .B(n25369), .C(n29228), .Y(n31361) );
  OAI21X1 U20857 ( .A(n23368), .B(n29262), .C(n21952), .Y(n31362) );
  OAI21X1 U20858 ( .A(n32355), .B(n29257), .C(n26334), .Y(n31363) );
  AOI21X1 U20859 ( .A(n26476), .B(n23367), .C(n24042), .Y(n31365) );
  NAND3X1 U20860 ( .A(n24073), .B(n24488), .C(n22806), .Y(n22201) );
  AOI22X1 U20861 ( .A(n29197), .B(n23367), .C(n25544), .D(n23368), .Y(n31372)
         );
  OAI21X1 U20862 ( .A(n31373), .B(n29239), .C(n23038), .Y(n31369) );
  NOR3X1 U20863 ( .A(n31368), .B(n29285), .C(n31369), .Y(n31370) );
  NAND3X1 U20864 ( .A(n21465), .B(n22449), .C(n31370), .Y(n22200) );
  AOI21X1 U20865 ( .A(n29317), .B(n26863), .C(n29279), .Y(n31379) );
  AOI22X1 U20866 ( .A(n25962), .B(n23367), .C(n25785), .D(n23368), .Y(n31378)
         );
  OAI21X1 U20867 ( .A(n25280), .B(n25758), .C(n23126), .Y(n31376) );
  NAND3X1 U20868 ( .A(n24208), .B(n24398), .C(n22852), .Y(n22199) );
  AOI22X1 U20869 ( .A(n26321), .B(n23370), .C(n26024), .D(n32359), .Y(n31387)
         );
  AOI21X1 U20870 ( .A(n29268), .B(n25370), .C(n20834), .Y(n31381) );
  OAI21X1 U20871 ( .A(n23370), .B(n29262), .C(n21953), .Y(n31382) );
  OAI21X1 U20872 ( .A(n32359), .B(n29257), .C(n26324), .Y(n31383) );
  AOI21X1 U20873 ( .A(n26475), .B(n23369), .C(n24043), .Y(n31385) );
  NAND3X1 U20874 ( .A(n24074), .B(n24489), .C(n22807), .Y(n22205) );
  AOI22X1 U20875 ( .A(n20997), .B(n23369), .C(n25567), .D(n23370), .Y(n31392)
         );
  OAI21X1 U20876 ( .A(n31393), .B(n29239), .C(n23039), .Y(n31389) );
  NOR3X1 U20877 ( .A(n31389), .B(n29285), .C(n31388), .Y(n31390) );
  NAND3X1 U20878 ( .A(n31390), .B(n21467), .C(n22452), .Y(n22204) );
  AOI21X1 U20879 ( .A(n29317), .B(n26807), .C(n29279), .Y(n31400) );
  AOI22X1 U20880 ( .A(n25961), .B(n23369), .C(n25787), .D(n23370), .Y(n31399)
         );
  OAI21X1 U20881 ( .A(n25282), .B(n29245), .C(n23136), .Y(n31396) );
  NAND3X1 U20882 ( .A(n24209), .B(n24400), .C(n22853), .Y(n22203) );
  AOI22X1 U20883 ( .A(n26314), .B(n23372), .C(n26026), .D(n32363), .Y(n31407)
         );
  AOI21X1 U20884 ( .A(n29267), .B(n25371), .C(n26290), .Y(n31401) );
  OAI21X1 U20885 ( .A(n23372), .B(n29262), .C(n21954), .Y(n31402) );
  OAI21X1 U20886 ( .A(n32363), .B(n29257), .C(n26326), .Y(n31403) );
  AOI21X1 U20887 ( .A(n26476), .B(n23371), .C(n22241), .Y(n31405) );
  NAND3X1 U20888 ( .A(n24075), .B(n24490), .C(n22808), .Y(n22209) );
  AOI22X1 U20889 ( .A(n20820), .B(n23371), .C(n25534), .D(n23372), .Y(n31412)
         );
  OAI21X1 U20890 ( .A(n31413), .B(n29239), .C(n23040), .Y(n31409) );
  NOR3X1 U20891 ( .A(n31409), .B(n29285), .C(n31408), .Y(n31410) );
  NAND3X1 U20892 ( .A(n31410), .B(n21469), .C(n22745), .Y(n22208) );
  AOI21X1 U20893 ( .A(n29317), .B(n26755), .C(n29279), .Y(n31420) );
  AOI22X1 U20894 ( .A(n25960), .B(n23371), .C(n25820), .D(n23372), .Y(n31419)
         );
  OAI21X1 U20895 ( .A(n25284), .B(n29246), .C(n23168), .Y(n31416) );
  NAND3X1 U20896 ( .A(n24210), .B(n24402), .C(n22854), .Y(n22207) );
  AOI22X1 U20897 ( .A(n26318), .B(n23374), .C(n26021), .D(n32367), .Y(n31428)
         );
  OAI21X1 U20898 ( .A(n23374), .B(n29262), .C(n31422), .Y(n31423) );
  OAI21X1 U20899 ( .A(n32367), .B(n29257), .C(n26327), .Y(n31424) );
  AOI21X1 U20900 ( .A(n26474), .B(n23373), .C(n22245), .Y(n31426) );
  NAND3X1 U20901 ( .A(n24076), .B(n24491), .C(n22809), .Y(n22213) );
  AOI22X1 U20902 ( .A(n20819), .B(n23373), .C(n25537), .D(n23374), .Y(n31433)
         );
  OAI21X1 U20903 ( .A(n31434), .B(n29239), .C(n23041), .Y(n31430) );
  NOR3X1 U20904 ( .A(n31430), .B(n29285), .C(n31429), .Y(n31431) );
  NAND3X1 U20905 ( .A(n31431), .B(n21472), .C(n22746), .Y(n22212) );
  AOI21X1 U20906 ( .A(n29317), .B(n26712), .C(n29279), .Y(n31441) );
  AOI22X1 U20907 ( .A(n25945), .B(n23373), .C(n25820), .D(n23374), .Y(n31440)
         );
  OAI21X1 U20908 ( .A(n25286), .B(n29245), .C(n23170), .Y(n31437) );
  NAND3X1 U20909 ( .A(n24211), .B(n24404), .C(n22855), .Y(n22211) );
  AOI22X1 U20910 ( .A(n26317), .B(n23376), .C(n25997), .D(n32371), .Y(n31448)
         );
  OAI21X1 U20911 ( .A(n23376), .B(n29262), .C(n31442), .Y(n31443) );
  OAI21X1 U20912 ( .A(n32371), .B(n29257), .C(n26331), .Y(n31444) );
  AOI21X1 U20913 ( .A(n26475), .B(n23375), .C(n22246), .Y(n31446) );
  NAND3X1 U20914 ( .A(n24078), .B(n24492), .C(n22810), .Y(n22217) );
  AOI22X1 U20915 ( .A(n20820), .B(n23375), .C(n25562), .D(n23376), .Y(n31452)
         );
  OAI21X1 U20916 ( .A(n31453), .B(n29239), .C(n23042), .Y(n31449) );
  NOR3X1 U20917 ( .A(n31455), .B(n29285), .C(n31449), .Y(n31450) );
  NAND3X1 U20918 ( .A(n21475), .B(n31450), .C(n22747), .Y(n22216) );
  AOI21X1 U20919 ( .A(n29317), .B(n26679), .C(n29279), .Y(n31459) );
  AOI22X1 U20920 ( .A(n25949), .B(n23375), .C(n25786), .D(n23376), .Y(n31458)
         );
  OAI21X1 U20921 ( .A(n25288), .B(n25758), .C(n23172), .Y(n31456) );
  NAND3X1 U20922 ( .A(n24212), .B(n24406), .C(n22856), .Y(n22215) );
  AOI22X1 U20923 ( .A(n26305), .B(n23378), .C(n25998), .D(n32375), .Y(n31467)
         );
  AOI21X1 U20924 ( .A(n29267), .B(n25374), .C(n29228), .Y(n31461) );
  OAI21X1 U20925 ( .A(n23378), .B(n29262), .C(n21955), .Y(n31462) );
  OAI21X1 U20926 ( .A(n32375), .B(n29257), .C(n26324), .Y(n31463) );
  AOI21X1 U20927 ( .A(n26479), .B(n23377), .C(n24044), .Y(n31465) );
  NAND3X1 U20928 ( .A(n22654), .B(n24493), .C(n24079), .Y(n22221) );
  AOI22X1 U20929 ( .A(n29233), .B(n23377), .C(n25566), .D(n23378), .Y(n31472)
         );
  OAI21X1 U20930 ( .A(n31473), .B(n29239), .C(n23043), .Y(n31469) );
  NOR3X1 U20931 ( .A(n31469), .B(n29285), .C(n31468), .Y(n31470) );
  NAND3X1 U20932 ( .A(n24081), .B(n21478), .C(n31470), .Y(n22220) );
  AOI21X1 U20933 ( .A(n29317), .B(n26647), .C(n29279), .Y(n31480) );
  AOI22X1 U20934 ( .A(n25955), .B(n23377), .C(n25818), .D(n23378), .Y(n31479)
         );
  OAI21X1 U20935 ( .A(n25289), .B(n29244), .C(n23138), .Y(n31476) );
  NAND3X1 U20936 ( .A(n24213), .B(n24408), .C(n22857), .Y(n22219) );
  AOI22X1 U20937 ( .A(n26305), .B(n23380), .C(n25999), .D(n32379), .Y(n31487)
         );
  AOI21X1 U20938 ( .A(n29267), .B(n25375), .C(n29194), .Y(n31481) );
  OAI21X1 U20939 ( .A(n23380), .B(n29262), .C(n21956), .Y(n31482) );
  OAI21X1 U20940 ( .A(n32379), .B(n29257), .C(n26330), .Y(n31483) );
  AOI21X1 U20941 ( .A(n26474), .B(n23379), .C(n23438), .Y(n31485) );
  NAND3X1 U20942 ( .A(n24083), .B(n24494), .C(n22811), .Y(n22225) );
  AOI22X1 U20943 ( .A(n29233), .B(n23379), .C(n25564), .D(n23380), .Y(n31491)
         );
  OAI21X1 U20944 ( .A(n31492), .B(n29239), .C(n25842), .Y(n31488) );
  NOR3X1 U20945 ( .A(n25843), .B(n29285), .C(n31488), .Y(n31489) );
  NAND3X1 U20946 ( .A(n24085), .B(n21481), .C(n31489), .Y(n22224) );
  AOI21X1 U20947 ( .A(n29317), .B(n26621), .C(n29279), .Y(n31498) );
  AOI22X1 U20948 ( .A(n25942), .B(n23379), .C(n25819), .D(n23380), .Y(n31497)
         );
  OAI21X1 U20949 ( .A(n25291), .B(n25757), .C(n22981), .Y(n31494) );
  NAND3X1 U20950 ( .A(n24214), .B(n24409), .C(n22858), .Y(n22223) );
  AOI22X1 U20951 ( .A(n26307), .B(n23383), .C(n26000), .D(n32383), .Y(n31505)
         );
  OAI21X1 U20952 ( .A(n23383), .B(n29262), .C(n31500), .Y(n31501) );
  OAI21X1 U20953 ( .A(n32383), .B(n29257), .C(n26327), .Y(n31502) );
  AOI21X1 U20954 ( .A(n26457), .B(n23382), .C(n25461), .Y(n31503) );
  AOI22X1 U20955 ( .A(n20826), .B(n23382), .C(n25563), .D(n23383), .Y(n31510)
         );
  OAI21X1 U20956 ( .A(n31511), .B(n29239), .C(n23116), .Y(n31507) );
  NOR3X1 U20957 ( .A(n29285), .B(n31506), .C(n31507), .Y(n31508) );
  NAND3X1 U20958 ( .A(n24087), .B(n21484), .C(n31508), .Y(n22228) );
  AOI21X1 U20959 ( .A(n29317), .B(n26596), .C(n29279), .Y(n31517) );
  AOI22X1 U20960 ( .A(n25954), .B(n23382), .C(n25818), .D(n23383), .Y(n31516)
         );
  OAI21X1 U20961 ( .A(n25293), .B(n29245), .C(n23115), .Y(n31514) );
  NAND3X1 U20962 ( .A(n24215), .B(n24411), .C(n22859), .Y(n22227) );
  AOI22X1 U20963 ( .A(n26314), .B(n23385), .C(n26029), .D(n32387), .Y(n31524)
         );
  AOI21X1 U20964 ( .A(n29267), .B(n25377), .C(n26280), .Y(n31518) );
  OAI21X1 U20965 ( .A(n23385), .B(n29262), .C(n21957), .Y(n31519) );
  OAI21X1 U20966 ( .A(n32387), .B(n29257), .C(n26323), .Y(n31520) );
  AOI21X1 U20967 ( .A(n26465), .B(n23384), .C(n22250), .Y(n31522) );
  NAND3X1 U20968 ( .A(n24089), .B(n23461), .C(n22812), .Y(n22233) );
  AOI22X1 U20969 ( .A(n21003), .B(n23384), .C(n25561), .D(n23385), .Y(n31529)
         );
  OAI21X1 U20970 ( .A(n31530), .B(n29240), .C(n23044), .Y(n31526) );
  NOR3X1 U20971 ( .A(n31525), .B(n29286), .C(n31526), .Y(n31527) );
  NAND3X1 U20972 ( .A(n24091), .B(n21393), .C(n31527), .Y(n22232) );
  AOI21X1 U20973 ( .A(n29317), .B(n27163), .C(n29279), .Y(n31536) );
  AOI22X1 U20974 ( .A(n25937), .B(n23384), .C(n25817), .D(n23385), .Y(n31535)
         );
  OAI21X1 U20975 ( .A(n25295), .B(n25758), .C(n23174), .Y(n31533) );
  NAND3X1 U20976 ( .A(n24216), .B(n24413), .C(n22860), .Y(n22231) );
  AOI22X1 U20977 ( .A(n26307), .B(n23387), .C(n25989), .D(n32391), .Y(n31544)
         );
  AOI21X1 U20978 ( .A(n29267), .B(n25378), .C(n21078), .Y(n31538) );
  OAI21X1 U20979 ( .A(n23387), .B(n29262), .C(n21958), .Y(n31539) );
  OAI21X1 U20980 ( .A(n32391), .B(n29257), .C(n26324), .Y(n31540) );
  AOI21X1 U20981 ( .A(n26467), .B(n23386), .C(n22254), .Y(n31542) );
  AOI22X1 U20982 ( .A(n20826), .B(n23386), .C(n25560), .D(n23387), .Y(n31549)
         );
  OAI21X1 U20983 ( .A(n31550), .B(n29240), .C(n23045), .Y(n31546) );
  NOR3X1 U20984 ( .A(n31546), .B(n29286), .C(n31545), .Y(n31547) );
  NAND3X1 U20985 ( .A(n24092), .B(n24495), .C(n31547), .Y(n22236) );
  AOI21X1 U20986 ( .A(n29318), .B(n27067), .C(n29279), .Y(n31557) );
  AOI22X1 U20987 ( .A(n25953), .B(n23386), .C(n25800), .D(n23387), .Y(n31556)
         );
  OAI21X1 U20988 ( .A(n25297), .B(n29246), .C(n23176), .Y(n31553) );
  NAND3X1 U20989 ( .A(n24217), .B(n24414), .C(n22861), .Y(n22235) );
  AOI22X1 U20990 ( .A(n26319), .B(n23389), .C(n25990), .D(n32395), .Y(n31564)
         );
  AOI21X1 U20991 ( .A(n29267), .B(n25379), .C(n20840), .Y(n31558) );
  OAI21X1 U20992 ( .A(n23389), .B(n29262), .C(n21959), .Y(n31559) );
  OAI21X1 U20993 ( .A(n32395), .B(n29257), .C(n26324), .Y(n31560) );
  AOI21X1 U20994 ( .A(n26467), .B(n23388), .C(n22258), .Y(n31562) );
  AOI22X1 U20995 ( .A(n21001), .B(n23388), .C(n25562), .D(n23389), .Y(n31569)
         );
  OAI21X1 U20996 ( .A(n31570), .B(n29240), .C(n23199), .Y(n31566) );
  NOR3X1 U20997 ( .A(n31565), .B(n29286), .C(n31566), .Y(n31567) );
  NAND3X1 U20998 ( .A(n24094), .B(n24496), .C(n31567), .Y(n22240) );
  AOI21X1 U20999 ( .A(n29318), .B(n26987), .C(n29279), .Y(n31577) );
  AOI22X1 U21000 ( .A(n25952), .B(n23388), .C(n25823), .D(n23389), .Y(n31576)
         );
  OAI21X1 U21001 ( .A(n25299), .B(n29245), .C(n23178), .Y(n31573) );
  NAND3X1 U21002 ( .A(n24218), .B(n24416), .C(n22862), .Y(n22239) );
  AOI22X1 U21003 ( .A(n26321), .B(n23391), .C(n25991), .D(n32399), .Y(n31585)
         );
  OAI21X1 U21004 ( .A(n23391), .B(n29262), .C(n31579), .Y(n31580) );
  OAI21X1 U21005 ( .A(n32399), .B(n29257), .C(n26324), .Y(n31581) );
  AOI21X1 U21006 ( .A(n26461), .B(n23390), .C(n23439), .Y(n31583) );
  AOI22X1 U21007 ( .A(n20829), .B(n23390), .C(n25559), .D(n23391), .Y(n31590)
         );
  OAI21X1 U21008 ( .A(n31591), .B(n29240), .C(n25182), .Y(n31587) );
  NOR3X1 U21009 ( .A(n31586), .B(n29286), .C(n31587), .Y(n31588) );
  NAND3X1 U21010 ( .A(n24096), .B(n24497), .C(n31588), .Y(n22244) );
  AOI21X1 U21011 ( .A(n29318), .B(n26922), .C(n29279), .Y(n31597) );
  AOI22X1 U21012 ( .A(n25943), .B(n23390), .C(n25824), .D(n23391), .Y(n31596)
         );
  OAI21X1 U21013 ( .A(n25301), .B(n25758), .C(n23127), .Y(n31594) );
  NAND3X1 U21014 ( .A(n24219), .B(n24418), .C(n22863), .Y(n22243) );
  AOI22X1 U21015 ( .A(n26322), .B(n23393), .C(n25992), .D(n32403), .Y(n31604)
         );
  AOI21X1 U21016 ( .A(n29267), .B(n25381), .C(n26298), .Y(n31599) );
  OAI21X1 U21017 ( .A(n23393), .B(n29263), .C(n21960), .Y(n31600) );
  OAI21X1 U21018 ( .A(n32403), .B(n29258), .C(n26324), .Y(n31601) );
  AOI21X1 U21019 ( .A(n26466), .B(n23392), .C(n25669), .Y(n31602) );
  NAND3X1 U21020 ( .A(n22455), .B(n23462), .C(n24852), .Y(n22249) );
  AOI22X1 U21021 ( .A(n20824), .B(n23392), .C(n25561), .D(n23393), .Y(n31609)
         );
  OAI21X1 U21022 ( .A(n31610), .B(n29240), .C(n23046), .Y(n31606) );
  NOR3X1 U21023 ( .A(n31605), .B(n29286), .C(n31606), .Y(n31607) );
  NAND3X1 U21024 ( .A(n24098), .B(n24498), .C(n31607), .Y(n22248) );
  AOI21X1 U21025 ( .A(n29318), .B(n26862), .C(n29279), .Y(n31617) );
  AOI22X1 U21026 ( .A(n25950), .B(n23392), .C(n25822), .D(n23393), .Y(n31616)
         );
  OAI21X1 U21027 ( .A(n25303), .B(n25856), .C(n25670), .Y(n31613) );
  NAND3X1 U21028 ( .A(n24220), .B(n24420), .C(n22864), .Y(n22247) );
  AOI22X1 U21029 ( .A(n26473), .B(n32407), .C(n26320), .D(n23395), .Y(n31623)
         );
  OAI21X1 U21030 ( .A(n23394), .B(n29258), .C(n26327), .Y(n31618) );
  AOI21X1 U21031 ( .A(n29267), .B(n25383), .C(n21056), .Y(n31619) );
  OAI21X1 U21032 ( .A(n23395), .B(n29263), .C(n21961), .Y(n31620) );
  NOR3X1 U21033 ( .A(n27226), .B(n31851), .C(n31625), .Y(n31621) );
  NAND3X1 U21034 ( .A(n31621), .B(n24499), .C(n22458), .Y(n22253) );
  AOI22X1 U21035 ( .A(n25542), .B(n23395), .C(n25902), .D(n23394), .Y(n31629)
         );
  NOR3X1 U21036 ( .A(n31626), .B(n29277), .C(n31625), .Y(n31627) );
  NAND3X1 U21037 ( .A(n24100), .B(n23463), .C(n31627), .Y(n22252) );
  AOI21X1 U21038 ( .A(n25949), .B(n32407), .C(n29287), .Y(n31634) );
  AOI22X1 U21039 ( .A(n25814), .B(n23395), .C(n25854), .D(n23394), .Y(n31633)
         );
  OAI21X1 U21040 ( .A(n31624), .B(n29210), .C(n23047), .Y(n31631) );
  NAND3X1 U21041 ( .A(n24221), .B(n24421), .C(n22865), .Y(n22251) );
  AOI22X1 U21042 ( .A(n26320), .B(n23397), .C(n25993), .D(n32411), .Y(n31641)
         );
  OAI21X1 U21043 ( .A(n23397), .B(n29263), .C(n31636), .Y(n31637) );
  OAI21X1 U21044 ( .A(n32411), .B(n29258), .C(n26324), .Y(n31638) );
  AOI21X1 U21045 ( .A(n26465), .B(n23396), .C(n25606), .Y(n31639) );
  NAND3X1 U21046 ( .A(n22461), .B(n24500), .C(n24854), .Y(n22257) );
  AOI22X1 U21047 ( .A(n21002), .B(n23396), .C(n25563), .D(n23397), .Y(n31645)
         );
  OAI21X1 U21048 ( .A(n31646), .B(n29240), .C(n23049), .Y(n31642) );
  NOR3X1 U21049 ( .A(n29286), .B(n21033), .C(n31642), .Y(n31643) );
  NAND3X1 U21050 ( .A(n31643), .B(n24501), .C(n24102), .Y(n22256) );
  AOI21X1 U21051 ( .A(n29318), .B(n26806), .C(n29279), .Y(n31653) );
  AOI22X1 U21052 ( .A(n25942), .B(n23396), .C(n25799), .D(n23397), .Y(n31652)
         );
  OAI21X1 U21053 ( .A(n25305), .B(n29246), .C(n25674), .Y(n31649) );
  NAND3X1 U21054 ( .A(n24222), .B(n24422), .C(n22866), .Y(n22255) );
  AOI22X1 U21055 ( .A(n26471), .B(n32415), .C(n26309), .D(n23399), .Y(n31659)
         );
  OAI21X1 U21056 ( .A(n23398), .B(n29258), .C(n26324), .Y(n31654) );
  AOI21X1 U21057 ( .A(n29266), .B(n27009), .C(n26302), .Y(n31655) );
  OAI21X1 U21058 ( .A(n23399), .B(n29263), .C(n21962), .Y(n31656) );
  NOR3X1 U21059 ( .A(n31661), .B(n31851), .C(n31662), .Y(n31657) );
  NAND3X1 U21060 ( .A(n31657), .B(n24502), .C(n22464), .Y(n22261) );
  AOI22X1 U21061 ( .A(n25543), .B(n23399), .C(n25925), .D(n23398), .Y(n31666)
         );
  OAI21X1 U21062 ( .A(n27009), .B(n29208), .C(n23050), .Y(n31663) );
  NOR3X1 U21063 ( .A(n29277), .B(n31662), .C(n31663), .Y(n31664) );
  NAND3X1 U21064 ( .A(n22467), .B(n24503), .C(n31664), .Y(n22260) );
  AOI21X1 U21065 ( .A(n25948), .B(n32415), .C(n29287), .Y(n31671) );
  AOI22X1 U21066 ( .A(n25813), .B(n23399), .C(n25854), .D(n23398), .Y(n31670)
         );
  OAI21X1 U21067 ( .A(n31660), .B(n29210), .C(n23052), .Y(n31668) );
  NAND3X1 U21068 ( .A(n24223), .B(n24423), .C(n22867), .Y(n22259) );
  AOI22X1 U21069 ( .A(n26317), .B(n23401), .C(n25994), .D(n32419), .Y(n31679)
         );
  AOI21X1 U21070 ( .A(n29266), .B(n25385), .C(n26291), .Y(n31673) );
  OAI21X1 U21071 ( .A(n23401), .B(n29263), .C(n21963), .Y(n31674) );
  OAI21X1 U21072 ( .A(n32419), .B(n29258), .C(n26336), .Y(n31675) );
  AOI21X1 U21073 ( .A(n20821), .B(n23400), .C(n22262), .Y(n31677) );
  AOI22X1 U21074 ( .A(n29232), .B(n23400), .C(n25559), .D(n23401), .Y(n31684)
         );
  OAI21X1 U21075 ( .A(n31685), .B(n29240), .C(n23053), .Y(n31681) );
  NOR3X1 U21076 ( .A(n31681), .B(n29286), .C(n31680), .Y(n31682) );
  NAND3X1 U21077 ( .A(n24104), .B(n24504), .C(n31682), .Y(n22264) );
  AOI21X1 U21078 ( .A(n29318), .B(n26754), .C(n29280), .Y(n31691) );
  AOI22X1 U21079 ( .A(n25941), .B(n23400), .C(n25796), .D(n23401), .Y(n31690)
         );
  OAI21X1 U21080 ( .A(n25307), .B(n25857), .C(n23180), .Y(n31688) );
  NAND3X1 U21081 ( .A(n24224), .B(n24425), .C(n22868), .Y(n22263) );
  AOI22X1 U21082 ( .A(n32423), .B(n26475), .C(n26318), .D(n23403), .Y(n31697)
         );
  OAI21X1 U21083 ( .A(n23402), .B(n29258), .C(n26328), .Y(n31692) );
  AOI21X1 U21084 ( .A(n29266), .B(n26944), .C(n26296), .Y(n31693) );
  OAI21X1 U21085 ( .A(n23403), .B(n29263), .C(n21964), .Y(n31694) );
  NOR3X1 U21086 ( .A(n31707), .B(n31897), .C(n31700), .Y(n31695) );
  NAND3X1 U21087 ( .A(n31695), .B(n24505), .C(n22470), .Y(n22269) );
  AOI22X1 U21088 ( .A(n25541), .B(n23403), .C(n25926), .D(n23402), .Y(n31704)
         );
  OAI21X1 U21089 ( .A(n26944), .B(n29208), .C(n23054), .Y(n31701) );
  NOR3X1 U21090 ( .A(n29277), .B(n31700), .C(n31701), .Y(n31702) );
  NAND3X1 U21091 ( .A(n22473), .B(n24506), .C(n31702), .Y(n22268) );
  AOI21X1 U21092 ( .A(n25952), .B(n32423), .C(n29287), .Y(n31710) );
  AOI22X1 U21093 ( .A(n25812), .B(n23403), .C(n25854), .D(n23402), .Y(n31709)
         );
  OAI21X1 U21094 ( .A(n31698), .B(n29210), .C(n23056), .Y(n31706) );
  NAND3X1 U21095 ( .A(n24225), .B(n24426), .C(n22869), .Y(n22267) );
  AOI22X1 U21096 ( .A(n26314), .B(n23405), .C(n25995), .D(n32427), .Y(n31718)
         );
  AOI21X1 U21097 ( .A(n29266), .B(n25386), .C(n26283), .Y(n31712) );
  OAI21X1 U21098 ( .A(n23405), .B(n29263), .C(n21965), .Y(n31713) );
  OAI21X1 U21099 ( .A(n32427), .B(n29258), .C(n26327), .Y(n31714) );
  AOI21X1 U21100 ( .A(n26453), .B(n23404), .C(n22265), .Y(n31716) );
  AOI22X1 U21101 ( .A(n20827), .B(n23404), .C(n25560), .D(n23405), .Y(n31723)
         );
  OAI21X1 U21102 ( .A(n31724), .B(n29240), .C(n22999), .Y(n31720) );
  NOR3X1 U21103 ( .A(n29286), .B(n31720), .C(n31719), .Y(n31721) );
  NAND3X1 U21104 ( .A(n24105), .B(n24507), .C(n31721), .Y(n22272) );
  AOI21X1 U21105 ( .A(n29318), .B(n26711), .C(n29280), .Y(n31731) );
  AOI22X1 U21106 ( .A(n25947), .B(n23404), .C(n25822), .D(n23405), .Y(n31730)
         );
  OAI21X1 U21107 ( .A(n25308), .B(n25757), .C(n23181), .Y(n31727) );
  NAND3X1 U21108 ( .A(n24226), .B(n24428), .C(n22870), .Y(n22271) );
  AOI22X1 U21109 ( .A(n26472), .B(n23407), .C(n26309), .D(n23408), .Y(n31737)
         );
  OAI21X1 U21110 ( .A(n23406), .B(n29258), .C(n26330), .Y(n31732) );
  AOI21X1 U21111 ( .A(n29266), .B(n25387), .C(n20834), .Y(n31733) );
  OAI21X1 U21112 ( .A(n23408), .B(n29263), .C(n21966), .Y(n31734) );
  NOR3X1 U21113 ( .A(n27227), .B(n31851), .C(n31739), .Y(n31735) );
  NAND3X1 U21114 ( .A(n31735), .B(n24508), .C(n22476), .Y(n22277) );
  AOI22X1 U21115 ( .A(n25558), .B(n23408), .C(n25927), .D(n23406), .Y(n31743)
         );
  NOR3X1 U21116 ( .A(n31739), .B(n29277), .C(n31740), .Y(n31741) );
  NAND3X1 U21117 ( .A(n24107), .B(n24509), .C(n31741), .Y(n22276) );
  AOI21X1 U21118 ( .A(n25940), .B(n23407), .C(n29287), .Y(n31748) );
  AOI22X1 U21119 ( .A(n25811), .B(n23408), .C(n25854), .D(n23406), .Y(n31747)
         );
  OAI21X1 U21120 ( .A(n31738), .B(n29210), .C(n23057), .Y(n31745) );
  NAND3X1 U21121 ( .A(n24227), .B(n24429), .C(n22871), .Y(n22275) );
  AOI22X1 U21122 ( .A(n26320), .B(n23410), .C(n26021), .D(n32434), .Y(n31756)
         );
  AOI21X1 U21123 ( .A(n29266), .B(n25388), .C(n20834), .Y(n31750) );
  OAI21X1 U21124 ( .A(n23410), .B(n29263), .C(n21967), .Y(n31751) );
  OAI21X1 U21125 ( .A(n32434), .B(n29258), .C(n26336), .Y(n31752) );
  AOI21X1 U21126 ( .A(n26454), .B(n23409), .C(n22266), .Y(n31754) );
  NAND3X1 U21127 ( .A(n24108), .B(n24510), .C(n22813), .Y(n22281) );
  AOI22X1 U21128 ( .A(n20825), .B(n23409), .C(n25550), .D(n23410), .Y(n31761)
         );
  OAI21X1 U21129 ( .A(n31762), .B(n29240), .C(n23059), .Y(n31758) );
  NOR3X1 U21130 ( .A(n31758), .B(n29286), .C(n31757), .Y(n31759) );
  NAND3X1 U21131 ( .A(n24109), .B(n22729), .C(n31759), .Y(n22280) );
  AOI21X1 U21132 ( .A(n29318), .B(n26678), .C(n29280), .Y(n31769) );
  AOI22X1 U21133 ( .A(n25939), .B(n23409), .C(n25792), .D(n23410), .Y(n31768)
         );
  OAI21X1 U21134 ( .A(n25310), .B(n29246), .C(n23183), .Y(n31765) );
  NAND3X1 U21135 ( .A(n24228), .B(n24431), .C(n22872), .Y(n22279) );
  AOI22X1 U21136 ( .A(n26449), .B(n32438), .C(n26308), .D(n23412), .Y(n31775)
         );
  OAI21X1 U21137 ( .A(n23411), .B(n29258), .C(n26328), .Y(n31770) );
  AOI21X1 U21138 ( .A(n29266), .B(n27104), .C(n26293), .Y(n31771) );
  OAI21X1 U21139 ( .A(n23412), .B(n29263), .C(n21968), .Y(n31772) );
  NOR3X1 U21140 ( .A(n31785), .B(n31897), .C(n31778), .Y(n31773) );
  NAND3X1 U21141 ( .A(n22479), .B(n24511), .C(n31773), .Y(n22285) );
  AOI22X1 U21142 ( .A(n25539), .B(n23412), .C(n25896), .D(n23411), .Y(n31782)
         );
  NAND3X1 U21143 ( .A(n22482), .B(n24512), .C(n21417), .Y(n22284) );
  AOI21X1 U21144 ( .A(n25945), .B(n32438), .C(n29287), .Y(n31788) );
  AOI22X1 U21145 ( .A(n25810), .B(n23412), .C(n25854), .D(n23411), .Y(n31787)
         );
  OAI21X1 U21146 ( .A(n31776), .B(n29210), .C(n23060), .Y(n31784) );
  NAND3X1 U21147 ( .A(n24229), .B(n24432), .C(n22873), .Y(n22283) );
  AOI22X1 U21148 ( .A(n26320), .B(n23414), .C(n26021), .D(n32442), .Y(n31796)
         );
  OAI21X1 U21149 ( .A(n23414), .B(n29263), .C(n31790), .Y(n31791) );
  OAI21X1 U21150 ( .A(n32442), .B(n29258), .C(n26336), .Y(n31792) );
  AOI21X1 U21151 ( .A(n26447), .B(n23413), .C(n24045), .Y(n31794) );
  NAND3X1 U21152 ( .A(n24110), .B(n24513), .C(n22814), .Y(n22289) );
  AOI22X1 U21153 ( .A(n29205), .B(n23413), .C(n25558), .D(n23414), .Y(n31801)
         );
  OAI21X1 U21154 ( .A(n31802), .B(n29240), .C(n23061), .Y(n31798) );
  NOR3X1 U21155 ( .A(n31797), .B(n29286), .C(n31798), .Y(n31799) );
  NAND3X1 U21156 ( .A(n24112), .B(n24514), .C(n31799), .Y(n22288) );
  AOI21X1 U21157 ( .A(n29318), .B(n26646), .C(n29280), .Y(n31808) );
  AOI22X1 U21158 ( .A(n25946), .B(n23413), .C(n25785), .D(n23414), .Y(n31807)
         );
  OAI21X1 U21159 ( .A(n25312), .B(n25857), .C(n23130), .Y(n31805) );
  NAND3X1 U21160 ( .A(n24230), .B(n24434), .C(n22874), .Y(n22287) );
  AOI22X1 U21161 ( .A(n26448), .B(n32446), .C(n26308), .D(n23416), .Y(n31814)
         );
  OAI21X1 U21162 ( .A(n23415), .B(n29258), .C(n26336), .Y(n31809) );
  AOI21X1 U21163 ( .A(n29266), .B(n26943), .C(n26287), .Y(n31810) );
  OAI21X1 U21164 ( .A(n23416), .B(n29263), .C(n21969), .Y(n31811) );
  NOR3X1 U21165 ( .A(n31824), .B(n31897), .C(n31817), .Y(n31812) );
  NAND3X1 U21166 ( .A(n31812), .B(n24515), .C(n22485), .Y(n22293) );
  AOI22X1 U21167 ( .A(n25539), .B(n23416), .C(n25928), .D(n23415), .Y(n31821)
         );
  OAI21X1 U21168 ( .A(n26943), .B(n29208), .C(n23062), .Y(n31818) );
  NOR3X1 U21169 ( .A(n29277), .B(n31817), .C(n31818), .Y(n31819) );
  NAND3X1 U21170 ( .A(n22488), .B(n24516), .C(n31819), .Y(n22292) );
  AOI21X1 U21171 ( .A(n25949), .B(n32446), .C(n29287), .Y(n31827) );
  AOI22X1 U21172 ( .A(n25805), .B(n23416), .C(n25854), .D(n23415), .Y(n31826)
         );
  OAI21X1 U21173 ( .A(n31815), .B(n29210), .C(n23064), .Y(n31823) );
  NAND3X1 U21174 ( .A(n24231), .B(n24435), .C(n22875), .Y(n22291) );
  AOI22X1 U21175 ( .A(n26322), .B(n23418), .C(n26020), .D(n32450), .Y(n31835)
         );
  AOI21X1 U21176 ( .A(n29266), .B(n25390), .C(n29194), .Y(n31829) );
  OAI21X1 U21177 ( .A(n23418), .B(n29261), .C(n21970), .Y(n31830) );
  OAI21X1 U21178 ( .A(n32450), .B(n29259), .C(n26329), .Y(n31831) );
  AOI21X1 U21179 ( .A(n26477), .B(n23417), .C(n24046), .Y(n31833) );
  NAND3X1 U21180 ( .A(n24113), .B(n24517), .C(n22815), .Y(n22297) );
  AOI22X1 U21181 ( .A(n29205), .B(n23417), .C(n25564), .D(n23418), .Y(n31840)
         );
  OAI21X1 U21182 ( .A(n31841), .B(n29240), .C(n23065), .Y(n31837) );
  NOR3X1 U21183 ( .A(n31836), .B(n29286), .C(n31837), .Y(n31838) );
  NAND3X1 U21184 ( .A(n24115), .B(n24518), .C(n31838), .Y(n22296) );
  AOI21X1 U21185 ( .A(n29318), .B(n26620), .C(n29280), .Y(n31847) );
  AOI22X1 U21186 ( .A(n25938), .B(n23417), .C(n25793), .D(n23418), .Y(n31846)
         );
  OAI21X1 U21187 ( .A(n25314), .B(n25857), .C(n23132), .Y(n31844) );
  NAND3X1 U21188 ( .A(n24232), .B(n24437), .C(n22876), .Y(n22295) );
  AOI22X1 U21189 ( .A(n23420), .B(n21004), .C(n26311), .D(n23421), .Y(n31854)
         );
  OAI21X1 U21190 ( .A(n23419), .B(n29259), .C(n26329), .Y(n31848) );
  OAI21X1 U21191 ( .A(n23421), .B(n29261), .C(n31849), .Y(n31850) );
  NOR3X1 U21192 ( .A(n27229), .B(n31851), .C(n31856), .Y(n31852) );
  NAND3X1 U21193 ( .A(n31852), .B(n24519), .C(n22491), .Y(n22301) );
  AOI22X1 U21194 ( .A(n25538), .B(n23421), .C(n25897), .D(n23419), .Y(n31860)
         );
  NOR3X1 U21195 ( .A(n31857), .B(n29277), .C(n31856), .Y(n31858) );
  NAND3X1 U21196 ( .A(n24117), .B(n24520), .C(n31858), .Y(n22300) );
  AOI21X1 U21197 ( .A(n25951), .B(n23420), .C(n29287), .Y(n31866) );
  AOI22X1 U21198 ( .A(n25804), .B(n23421), .C(n29247), .D(n23419), .Y(n31865)
         );
  OAI21X1 U21199 ( .A(n31855), .B(n29210), .C(n23066), .Y(n31863) );
  NAND3X1 U21200 ( .A(n24233), .B(n24438), .C(n22877), .Y(n22299) );
  AOI22X1 U21201 ( .A(n26314), .B(n23423), .C(n26033), .D(n32457), .Y(n31875)
         );
  OAI21X1 U21202 ( .A(n23423), .B(n29261), .C(n31869), .Y(n31870) );
  OAI21X1 U21203 ( .A(n32457), .B(n29259), .C(n26323), .Y(n31871) );
  AOI21X1 U21204 ( .A(n26472), .B(n23422), .C(n22270), .Y(n31873) );
  NAND3X1 U21205 ( .A(n24119), .B(n24521), .C(n22816), .Y(n22305) );
  AOI22X1 U21206 ( .A(n29205), .B(n23422), .C(n25566), .D(n23423), .Y(n31881)
         );
  OAI21X1 U21207 ( .A(n31882), .B(n29240), .C(n23210), .Y(n31878) );
  NOR3X1 U21208 ( .A(n29286), .B(n31878), .C(n31877), .Y(n31879) );
  NAND3X1 U21209 ( .A(n24121), .B(n24522), .C(n31879), .Y(n22304) );
  AOI21X1 U21210 ( .A(n29318), .B(n26595), .C(n29280), .Y(n31889) );
  AOI22X1 U21211 ( .A(n25940), .B(n23422), .C(n25792), .D(n23423), .Y(n31888)
         );
  OAI21X1 U21212 ( .A(n25316), .B(n25857), .C(n23185), .Y(n31886) );
  NAND3X1 U21213 ( .A(n24234), .B(n24440), .C(n22878), .Y(n22303) );
  AOI22X1 U21214 ( .A(n26320), .B(n34495), .C(n26015), .D(n32463), .Y(n31898)
         );
  OAI21X1 U21215 ( .A(n32463), .B(n29259), .C(n26334), .Y(n31893) );
  AOI22X1 U21216 ( .A(n29266), .B(n25433), .C(n29264), .D(n25397), .Y(n31895)
         );
  NAND3X1 U21217 ( .A(n22494), .B(n25129), .C(n31909), .Y(n22309) );
  AOI22X1 U21218 ( .A(n25541), .B(n34495), .C(n25895), .D(n32463), .Y(n31906)
         );
  OAI21X1 U21219 ( .A(n25434), .B(n29208), .C(n23087), .Y(n31903) );
  NOR3X1 U21220 ( .A(n31902), .B(n29277), .C(n31903), .Y(n31904) );
  NAND3X1 U21221 ( .A(n22497), .B(n24523), .C(n31904), .Y(n22308) );
  AOI22X1 U21222 ( .A(n34496), .B(n25944), .C(n34495), .D(n25798), .Y(n31911)
         );
  AOI22X1 U21223 ( .A(n25854), .B(n32463), .C(n29277), .D(n27179), .Y(n31910)
         );
  AOI22X1 U21224 ( .A(net96340), .B(n22794), .C(n29374), .D(n31912), .Y(n31915) );
  OR2X2 U21225 ( .A(n22102), .B(n27157), .Y(n31921) );
  AOI21X1 U21226 ( .A(n32101), .B(n27170), .C(n20815), .Y(n31920) );
  AOI22X1 U21227 ( .A(n29311), .B(n25007), .C(n29304), .D(n31917), .Y(n31918)
         );
  NAND3X1 U21228 ( .A(n22655), .B(n24524), .C(n24713), .Y(n22056) );
  AOI22X1 U21229 ( .A(n29311), .B(n25008), .C(n29304), .D(n25227), .Y(n31925)
         );
  NAND3X1 U21230 ( .A(n20996), .B(n24525), .C(n24714), .Y(n34507) );
  AOI21X1 U21231 ( .A(n32101), .B(n26861), .C(n32099), .Y(n31932) );
  AOI22X1 U21232 ( .A(n29311), .B(n25009), .C(n29304), .D(n25229), .Y(n31930)
         );
  NAND3X1 U21233 ( .A(n22656), .B(n24526), .C(n24715), .Y(n22066) );
  AOI22X1 U21234 ( .A(n29311), .B(n25010), .C(n29304), .D(n25231), .Y(n31935)
         );
  NAND3X1 U21235 ( .A(n20996), .B(n24527), .C(n24716), .Y(n34508) );
  AOI21X1 U21236 ( .A(n32101), .B(n26993), .C(n20816), .Y(n31942) );
  AOI22X1 U21237 ( .A(n29311), .B(n25011), .C(n29303), .D(n25233), .Y(n31940)
         );
  NAND3X1 U21238 ( .A(n24717), .B(n24528), .C(n22657), .Y(n22074) );
  AOI22X1 U21239 ( .A(n29311), .B(n25012), .C(n29303), .D(n25235), .Y(n31945)
         );
  NAND3X1 U21240 ( .A(n20996), .B(n24529), .C(n24718), .Y(n34509) );
  AOI21X1 U21241 ( .A(n32101), .B(n27073), .C(n20815), .Y(n31952) );
  AOI22X1 U21242 ( .A(n29311), .B(n25013), .C(n29303), .D(n25237), .Y(n31950)
         );
  NAND3X1 U21243 ( .A(n22658), .B(n24530), .C(n24719), .Y(n22082) );
  AOI22X1 U21244 ( .A(n29311), .B(n25014), .C(n29303), .D(n25239), .Y(n31956)
         );
  NAND3X1 U21245 ( .A(n20996), .B(n24531), .C(n24720), .Y(n34510) );
  AOI21X1 U21246 ( .A(n32101), .B(n27072), .C(n20981), .Y(n31963) );
  AOI22X1 U21247 ( .A(n29311), .B(n25015), .C(n29303), .D(n25241), .Y(n31961)
         );
  NAND3X1 U21248 ( .A(n22659), .B(n24532), .C(n24721), .Y(n22090) );
  AOI22X1 U21249 ( .A(n29311), .B(n25016), .C(n29303), .D(n25243), .Y(n31966)
         );
  NAND3X1 U21250 ( .A(n20990), .B(n24533), .C(n24722), .Y(n34511) );
  AOI21X1 U21251 ( .A(n32101), .B(n27169), .C(n20823), .Y(n31973) );
  AOI22X1 U21252 ( .A(n29311), .B(n25017), .C(n29303), .D(n25245), .Y(n31971)
         );
  NAND3X1 U21253 ( .A(n22660), .B(n24534), .C(n24723), .Y(n22098) );
  AOI22X1 U21254 ( .A(n29311), .B(n25018), .C(n29303), .D(n25247), .Y(n31975)
         );
  NAND3X1 U21255 ( .A(n20996), .B(n24535), .C(n24724), .Y(n34512) );
  AOI21X1 U21256 ( .A(n32101), .B(n26921), .C(n20816), .Y(n31982) );
  AOI22X1 U21257 ( .A(n29310), .B(n25019), .C(n29303), .D(n25249), .Y(n31980)
         );
  NAND3X1 U21258 ( .A(n22661), .B(n24536), .C(n24725), .Y(n22106) );
  AOI22X1 U21259 ( .A(n29310), .B(n25020), .C(n29303), .D(n25251), .Y(n31985)
         );
  NAND3X1 U21260 ( .A(n20989), .B(n24537), .C(n24726), .Y(n34513) );
  AOI21X1 U21261 ( .A(n32101), .B(n26992), .C(n20980), .Y(n31993) );
  AOI22X1 U21262 ( .A(n29310), .B(n25164), .C(n29303), .D(n25253), .Y(n31991)
         );
  NAND3X1 U21263 ( .A(n22662), .B(n24538), .C(n24727), .Y(n22114) );
  AOI22X1 U21264 ( .A(n29310), .B(n25021), .C(n29303), .D(n25255), .Y(n31996)
         );
  NAND3X1 U21265 ( .A(n20996), .B(n24539), .C(n24728), .Y(n34514) );
  AOI22X1 U21266 ( .A(n29310), .B(n25022), .C(n29302), .D(n25257), .Y(n31998)
         );
  NAND3X1 U21267 ( .A(n25741), .B(n24540), .C(n24729), .Y(n34515) );
  AOI22X1 U21268 ( .A(n29310), .B(n25023), .C(n29302), .D(n25085), .Y(n32001)
         );
  NAND3X1 U21269 ( .A(n25740), .B(n24541), .C(n24730), .Y(n34516) );
  AOI22X1 U21270 ( .A(n29310), .B(n25024), .C(n29302), .D(n25259), .Y(n32003)
         );
  NAND3X1 U21271 ( .A(n25735), .B(n24542), .C(n24731), .Y(n34517) );
  AOI22X1 U21272 ( .A(n29310), .B(n25025), .C(n25086), .D(n29302), .Y(n32006)
         );
  NAND3X1 U21273 ( .A(n25736), .B(n24543), .C(n24732), .Y(n34518) );
  AOI22X1 U21274 ( .A(n29310), .B(n25026), .C(n29302), .D(n25260), .Y(n32009)
         );
  NAND3X1 U21275 ( .A(n20983), .B(n24544), .C(n24733), .Y(n34519) );
  AOI22X1 U21276 ( .A(n29310), .B(n25027), .C(n25087), .D(n29302), .Y(n32012)
         );
  NAND3X1 U21277 ( .A(n25739), .B(n24545), .C(n24734), .Y(n34520) );
  AOI22X1 U21278 ( .A(n29310), .B(n25028), .C(n29302), .D(n25262), .Y(n32015)
         );
  NAND3X1 U21279 ( .A(n25737), .B(n24546), .C(n24735), .Y(n34521) );
  AOI22X1 U21280 ( .A(n29310), .B(n25029), .C(n25088), .D(n29302), .Y(n32018)
         );
  NAND3X1 U21281 ( .A(n25738), .B(n24547), .C(n24736), .Y(n34522) );
  AOI22X1 U21282 ( .A(n29310), .B(n25030), .C(n29302), .D(n25264), .Y(n32021)
         );
  NAND3X1 U21283 ( .A(n20996), .B(n24548), .C(n24737), .Y(n34523) );
  AOI22X1 U21284 ( .A(n29309), .B(n25165), .C(n29302), .D(n25089), .Y(n32024)
         );
  NAND3X1 U21285 ( .A(n20990), .B(n24549), .C(n24738), .Y(n34524) );
  AOI22X1 U21286 ( .A(n29309), .B(n25031), .C(n29302), .D(n25266), .Y(n32027)
         );
  NAND3X1 U21287 ( .A(n25742), .B(n24550), .C(n24739), .Y(n34525) );
  AOI22X1 U21288 ( .A(n29309), .B(n25032), .C(n25090), .D(n29302), .Y(n32030)
         );
  NAND3X1 U21289 ( .A(n25735), .B(n24551), .C(n24740), .Y(n34526) );
  AOI22X1 U21290 ( .A(n29309), .B(n25033), .C(n29301), .D(n25268), .Y(n32033)
         );
  NAND3X1 U21291 ( .A(n20990), .B(n24552), .C(n24741), .Y(n34527) );
  AOI22X1 U21292 ( .A(n29309), .B(n25034), .C(n29301), .D(n25091), .Y(n32036)
         );
  NAND3X1 U21293 ( .A(n20822), .B(n24553), .C(n24742), .Y(n34528) );
  AOI22X1 U21294 ( .A(n29309), .B(n25035), .C(n29301), .D(n25270), .Y(n32039)
         );
  NAND3X1 U21295 ( .A(n25735), .B(n24554), .C(n24743), .Y(n34529) );
  AOI22X1 U21296 ( .A(n29309), .B(n25036), .C(n29301), .D(n25205), .Y(n32043)
         );
  NAND3X1 U21297 ( .A(n25740), .B(n24555), .C(n24744), .Y(n34530) );
  AOI21X1 U21298 ( .A(n32101), .B(n26860), .C(n20981), .Y(n32049) );
  AOI22X1 U21299 ( .A(n29309), .B(n25037), .C(n29301), .D(n25272), .Y(n32047)
         );
  NAND3X1 U21300 ( .A(n22663), .B(n24556), .C(n24745), .Y(n22186) );
  AOI22X1 U21301 ( .A(n29309), .B(n25038), .C(n29301), .D(n25274), .Y(n32051)
         );
  NAND3X1 U21302 ( .A(n25740), .B(n24557), .C(n24746), .Y(n34531) );
  AOI21X1 U21303 ( .A(n32101), .B(n27071), .C(n20980), .Y(n32057) );
  AOI22X1 U21304 ( .A(n29309), .B(n25039), .C(n29301), .D(n25276), .Y(n32055)
         );
  NAND3X1 U21305 ( .A(n22664), .B(n24558), .C(n24747), .Y(n22194) );
  AOI22X1 U21306 ( .A(n29309), .B(n25040), .C(n29301), .D(n25278), .Y(n32058)
         );
  NAND3X1 U21307 ( .A(n25740), .B(n24559), .C(n24748), .Y(n34532) );
  AOI21X1 U21308 ( .A(n32101), .B(n27168), .C(n20987), .Y(n32064) );
  AOI22X1 U21309 ( .A(n29309), .B(n25041), .C(n29301), .D(n25280), .Y(n32062)
         );
  NAND3X1 U21310 ( .A(n22665), .B(n24560), .C(n24749), .Y(n22202) );
  AOI22X1 U21311 ( .A(n29309), .B(n25042), .C(n29301), .D(n25282), .Y(n32066)
         );
  NAND3X1 U21312 ( .A(n25736), .B(n24561), .C(n24750), .Y(n34533) );
  AOI21X1 U21313 ( .A(n32101), .B(n26927), .C(n20817), .Y(n32072) );
  AOI22X1 U21314 ( .A(n29308), .B(n25043), .C(n29301), .D(n25284), .Y(n32070)
         );
  NAND3X1 U21315 ( .A(n22666), .B(n24562), .C(n24751), .Y(n22210) );
  AOI22X1 U21316 ( .A(n29308), .B(n25044), .C(n29301), .D(n25286), .Y(n32074)
         );
  NAND3X1 U21317 ( .A(n25740), .B(n24563), .C(n24752), .Y(n34534) );
  AOI21X1 U21318 ( .A(n32101), .B(n26991), .C(n20817), .Y(n32080) );
  AOI22X1 U21319 ( .A(n29308), .B(n25045), .C(n29300), .D(n25288), .Y(n32078)
         );
  NAND3X1 U21320 ( .A(n22667), .B(n24564), .C(n24753), .Y(n22218) );
  AOI22X1 U21321 ( .A(n29308), .B(n25046), .C(n29300), .D(n25289), .Y(n32082)
         );
  NAND3X1 U21322 ( .A(n20985), .B(n24565), .C(n24754), .Y(n34535) );
  AOI21X1 U21323 ( .A(n32101), .B(n26926), .C(n32099), .Y(n32088) );
  AOI22X1 U21324 ( .A(n29308), .B(n25047), .C(n29300), .D(n25291), .Y(n32086)
         );
  NAND3X1 U21325 ( .A(n22668), .B(n24566), .C(n24755), .Y(n22226) );
  AOI22X1 U21326 ( .A(n29308), .B(n25048), .C(n29300), .D(n25293), .Y(n32089)
         );
  NAND3X1 U21327 ( .A(n20984), .B(n24567), .C(n24756), .Y(n34536) );
  AOI21X1 U21328 ( .A(n32101), .B(n27066), .C(n20823), .Y(n32095) );
  AOI22X1 U21329 ( .A(n29308), .B(n25049), .C(n29300), .D(n25295), .Y(n32093)
         );
  NAND3X1 U21330 ( .A(n22669), .B(n24568), .C(n24757), .Y(n22234) );
  AOI22X1 U21331 ( .A(n29308), .B(n25050), .C(n29300), .D(n25297), .Y(n32097)
         );
  NAND3X1 U21332 ( .A(n25740), .B(n24569), .C(n24758), .Y(n34537) );
  AOI21X1 U21333 ( .A(n32101), .B(n27167), .C(n20987), .Y(n32105) );
  AOI22X1 U21334 ( .A(n29308), .B(n25051), .C(n29300), .D(n25299), .Y(n32103)
         );
  NAND3X1 U21335 ( .A(n22670), .B(n24570), .C(n24759), .Y(n22242) );
  AOI22X1 U21336 ( .A(n29308), .B(n25052), .C(n29300), .D(n25301), .Y(n32107)
         );
  NAND3X1 U21337 ( .A(n25737), .B(n24571), .C(n24760), .Y(n34538) );
  AOI22X1 U21338 ( .A(n29308), .B(n25053), .C(n29300), .D(n25303), .Y(n32110)
         );
  NAND3X1 U21339 ( .A(n20986), .B(n24572), .C(n24761), .Y(n34539) );
  AOI22X1 U21340 ( .A(n29308), .B(n25054), .C(n29300), .D(n25092), .Y(n32113)
         );
  NAND3X1 U21341 ( .A(n25740), .B(n24573), .C(n24762), .Y(n34540) );
  AOI22X1 U21342 ( .A(n29308), .B(n25055), .C(n29300), .D(n25305), .Y(n32116)
         );
  NAND3X1 U21343 ( .A(n20989), .B(n24574), .C(n24763), .Y(n34541) );
  AOI22X1 U21344 ( .A(n29307), .B(n25056), .C(n25093), .D(n29300), .Y(n32119)
         );
  NAND3X1 U21345 ( .A(n20996), .B(n24575), .C(n24764), .Y(n34542) );
  AOI22X1 U21346 ( .A(n29307), .B(n25057), .C(n29299), .D(n25307), .Y(n32122)
         );
  NAND3X1 U21347 ( .A(n25739), .B(n24576), .C(n24765), .Y(n34543) );
  AOI22X1 U21348 ( .A(n29307), .B(n25058), .C(n29299), .D(n25094), .Y(n32125)
         );
  NAND3X1 U21349 ( .A(n25742), .B(n24577), .C(n24766), .Y(n34544) );
  AOI22X1 U21350 ( .A(n29307), .B(n25059), .C(n29299), .D(n25308), .Y(n32128)
         );
  NAND3X1 U21351 ( .A(n25738), .B(n24578), .C(n24767), .Y(n34545) );
  AOI22X1 U21352 ( .A(n29307), .B(n25060), .C(n29299), .D(n25095), .Y(n32130)
         );
  NAND3X1 U21353 ( .A(n20822), .B(n24579), .C(n24768), .Y(n34546) );
  AOI22X1 U21354 ( .A(n29307), .B(n25061), .C(n29299), .D(n25310), .Y(n32133)
         );
  NAND3X1 U21355 ( .A(n25740), .B(n24580), .C(n24769), .Y(n34547) );
  AOI22X1 U21356 ( .A(n29307), .B(n25062), .C(n29299), .D(n25096), .Y(n32136)
         );
  NAND3X1 U21357 ( .A(n20984), .B(n24581), .C(n24770), .Y(n34548) );
  AOI22X1 U21358 ( .A(n29307), .B(n25063), .C(n29299), .D(n25312), .Y(n32139)
         );
  NAND3X1 U21359 ( .A(n20985), .B(n24582), .C(n24771), .Y(n34549) );
  AOI22X1 U21360 ( .A(n29307), .B(n25064), .C(n29299), .D(n25097), .Y(n32142)
         );
  NAND3X1 U21361 ( .A(n20983), .B(n24583), .C(n24772), .Y(n34550) );
  AOI22X1 U21362 ( .A(n29307), .B(n25065), .C(n29299), .D(n25314), .Y(n32145)
         );
  NAND3X1 U21363 ( .A(n20996), .B(n24584), .C(n24773), .Y(n34551) );
  AOI22X1 U21364 ( .A(n29307), .B(n25066), .C(n29299), .D(n25098), .Y(n32147)
         );
  NAND3X1 U21365 ( .A(n25741), .B(n24585), .C(n24774), .Y(n34552) );
  AOI22X1 U21366 ( .A(n29307), .B(n25067), .C(n29299), .D(n25316), .Y(n32150)
         );
  NAND3X1 U21367 ( .A(n20986), .B(n24586), .C(n24775), .Y(n34553) );
  AOI22X1 U21368 ( .A(n29307), .B(n25398), .C(n29299), .D(n25449), .Y(n32155)
         );
  NAND3X1 U21369 ( .A(n25738), .B(n24587), .C(n24776), .Y(n34554) );
  AOI22X1 U21370 ( .A(T[5]), .B(n34613), .C(n23281), .D(n2256), .Y(n32158) );
  OAI21X1 U21371 ( .A(n27118), .B(n32159), .C(n21567), .Y(n32160) );
  AOI22X1 U21372 ( .A(n32157), .B(n32160), .C(n23425), .D(n27211), .Y(n32162)
         );
  AOI22X1 U21373 ( .A(n27263), .B(net124030), .C(n23276), .D(n26482), .Y(
        n32161) );
  AOI22X1 U21374 ( .A(T[4]), .B(n34613), .C(n23281), .D(n2255), .Y(n32163) );
  OAI21X1 U21375 ( .A(n27118), .B(n32164), .C(n21568), .Y(n32165) );
  AOI22X1 U21376 ( .A(n32157), .B(n32165), .C(n23425), .D(n25451), .Y(n32167)
         );
  AOI22X1 U21377 ( .A(n27263), .B(net104479), .C(n23276), .D(n2249), .Y(n32166) );
  AOI22X1 U21378 ( .A(T[3]), .B(n34613), .C(n23281), .D(n2254), .Y(n32168) );
  OAI21X1 U21379 ( .A(n27118), .B(n32169), .C(n21569), .Y(n32170) );
  AOI22X1 U21380 ( .A(n32157), .B(n32170), .C(n23425), .D(n28606), .Y(n32172)
         );
  AOI22X1 U21381 ( .A(n27263), .B(n28220), .C(n23276), .D(n27214), .Y(n32171)
         );
  AOI22X1 U21382 ( .A(T[2]), .B(n34613), .C(n23281), .D(n29185), .Y(n32173) );
  OAI21X1 U21383 ( .A(n27118), .B(n32174), .C(n21570), .Y(n32175) );
  AOI22X1 U21384 ( .A(n32157), .B(n32175), .C(n23425), .D(n28604), .Y(n32177)
         );
  AOI22X1 U21385 ( .A(n27263), .B(net149936), .C(n23276), .D(n26541), .Y(
        n32176) );
  AOI22X1 U21386 ( .A(T[1]), .B(n34613), .C(n23281), .D(n29182), .Y(n32178) );
  OAI21X1 U21387 ( .A(n27118), .B(n32179), .C(n21571), .Y(n32180) );
  AOI22X1 U21388 ( .A(n32157), .B(n32180), .C(n23425), .D(n26509), .Y(n32182)
         );
  AOI22X1 U21389 ( .A(n27263), .B(net105815), .C(n23276), .D(n26444), .Y(
        n32181) );
  AOI22X1 U21390 ( .A(T[0]), .B(n34613), .C(n23281), .D(alt5_net95652), .Y(
        n32183) );
  OAI21X1 U21391 ( .A(n27118), .B(n32184), .C(n21572), .Y(n32186) );
  AOI21X1 U21392 ( .A(n32157), .B(n32186), .C(n29318), .Y(n32189) );
  AOI22X1 U21393 ( .A(n27263), .B(net150130), .C(n23276), .D(n26174), .Y(
        n32187) );
  NAND3X1 U21394 ( .A(n24235), .B(n24588), .C(n24777), .Y(n21313) );
  NAND2X1 U21395 ( .A(n15195), .B(n32190), .Y(n22429) );
  OAI21X1 U21396 ( .A(n25003), .B(n25078), .C(n21991), .Y(n21852) );
  NAND2X1 U21397 ( .A(n29321), .B(n14097), .Y(n32193) );
  AOI21X1 U21398 ( .A(n31916), .B(n29323), .C(n14218), .Y(n32196) );
  NAND2X1 U21399 ( .A(n23311), .B(n14368), .Y(n32195) );
  AOI22X1 U21400 ( .A(n23310), .B(n14369), .C(n14371), .D(n25715), .Y(n32194)
         );
  NAND3X1 U21401 ( .A(n32196), .B(n32195), .C(n32194), .Y(n22436) );
  NAND3X1 U21402 ( .A(n25346), .B(n22730), .C(n29319), .Y(n22058) );
  AOI21X1 U21403 ( .A(n30670), .B(n29323), .C(n14218), .Y(n32203) );
  NAND2X1 U21404 ( .A(n32199), .B(n14371), .Y(n32202) );
  AOI22X1 U21405 ( .A(n23312), .B(n14368), .C(n32200), .D(n14369), .Y(n32201)
         );
  NAND3X1 U21406 ( .A(n32203), .B(n32202), .C(n32201), .Y(n22439) );
  AOI21X1 U21407 ( .A(n31927), .B(n29323), .C(n14218), .Y(n32208) );
  NAND2X1 U21408 ( .A(n32204), .B(n14371), .Y(n32207) );
  AOI22X1 U21409 ( .A(n23313), .B(n14368), .C(n32205), .D(n14369), .Y(n32206)
         );
  NAND3X1 U21410 ( .A(n32208), .B(n32207), .C(n32206), .Y(n22442) );
  AOI21X1 U21411 ( .A(n30713), .B(n29323), .C(n14218), .Y(n32213) );
  NAND2X1 U21412 ( .A(n32209), .B(n14371), .Y(n32212) );
  AOI22X1 U21413 ( .A(n23314), .B(n14368), .C(n32210), .D(n14369), .Y(n32211)
         );
  NAND3X1 U21414 ( .A(n32213), .B(n32212), .C(n32211), .Y(n22445) );
  AOI21X1 U21415 ( .A(n31937), .B(n29323), .C(n14218), .Y(n32218) );
  NAND2X1 U21416 ( .A(n32214), .B(n14371), .Y(n32217) );
  AOI22X1 U21417 ( .A(n23315), .B(n14368), .C(n32215), .D(n14369), .Y(n32216)
         );
  NAND3X1 U21418 ( .A(n32218), .B(n32217), .C(n32216), .Y(n22448) );
  AOI21X1 U21419 ( .A(n30753), .B(n29323), .C(n14218), .Y(n32223) );
  NAND2X1 U21420 ( .A(n32219), .B(n14371), .Y(n32222) );
  AOI22X1 U21421 ( .A(n23316), .B(n14368), .C(n32220), .D(n14369), .Y(n32221)
         );
  NAND3X1 U21422 ( .A(n32223), .B(n32222), .C(n32221), .Y(n22451) );
  AOI21X1 U21423 ( .A(n31947), .B(n29323), .C(n14218), .Y(n32228) );
  NAND2X1 U21424 ( .A(n32224), .B(n14371), .Y(n32227) );
  AOI22X1 U21425 ( .A(n23317), .B(n14368), .C(n32225), .D(n14369), .Y(n32226)
         );
  NAND3X1 U21426 ( .A(n32228), .B(n32227), .C(n32226), .Y(n22454) );
  AOI21X1 U21427 ( .A(n30793), .B(n29323), .C(n14218), .Y(n32233) );
  NAND2X1 U21428 ( .A(n32229), .B(n14371), .Y(n32232) );
  AOI22X1 U21429 ( .A(n31955), .B(n14368), .C(n32230), .D(n14369), .Y(n32231)
         );
  NAND3X1 U21430 ( .A(n32233), .B(n32232), .C(n32231), .Y(n22457) );
  AOI21X1 U21431 ( .A(n31958), .B(n29323), .C(n14218), .Y(n32238) );
  NAND2X1 U21432 ( .A(n32234), .B(n14371), .Y(n32237) );
  AOI22X1 U21433 ( .A(n23318), .B(n14368), .C(n32235), .D(n14369), .Y(n32236)
         );
  NAND3X1 U21434 ( .A(n32238), .B(n32237), .C(n32236), .Y(n22460) );
  AOI21X1 U21435 ( .A(n30833), .B(n29323), .C(n14218), .Y(n32243) );
  NAND2X1 U21436 ( .A(n32239), .B(n14371), .Y(n32242) );
  AOI22X1 U21437 ( .A(n23319), .B(n14368), .C(n32240), .D(n14369), .Y(n32241)
         );
  NAND3X1 U21438 ( .A(n32243), .B(n32242), .C(n32241), .Y(n22463) );
  AOI21X1 U21439 ( .A(n31968), .B(n29323), .C(n14218), .Y(n32248) );
  NAND2X1 U21440 ( .A(n32244), .B(n14371), .Y(n32247) );
  AOI22X1 U21441 ( .A(n23320), .B(n14368), .C(n32245), .D(n14369), .Y(n32246)
         );
  NAND3X1 U21442 ( .A(n32248), .B(n32247), .C(n32246), .Y(n22466) );
  AOI21X1 U21443 ( .A(n30873), .B(n29323), .C(n14218), .Y(n32253) );
  NAND2X1 U21444 ( .A(n32249), .B(n14371), .Y(n32252) );
  AOI22X1 U21445 ( .A(n23322), .B(n14368), .C(n32250), .D(n14369), .Y(n32251)
         );
  NAND3X1 U21446 ( .A(n32253), .B(n32252), .C(n32251), .Y(n22469) );
  AOI21X1 U21447 ( .A(n31977), .B(n29323), .C(n14218), .Y(n32258) );
  NAND2X1 U21448 ( .A(n32254), .B(n14371), .Y(n32257) );
  AOI22X1 U21449 ( .A(n23323), .B(n14368), .C(n32255), .D(n14369), .Y(n32256)
         );
  NAND3X1 U21450 ( .A(n32258), .B(n32257), .C(n32256), .Y(n22472) );
  AOI21X1 U21451 ( .A(n30914), .B(n29324), .C(n14218), .Y(n32263) );
  NAND2X1 U21452 ( .A(n32259), .B(n14371), .Y(n32262) );
  AOI22X1 U21453 ( .A(n23324), .B(n14368), .C(n32260), .D(n14369), .Y(n32261)
         );
  NAND3X1 U21454 ( .A(n32263), .B(n32262), .C(n32261), .Y(n22475) );
  AOI21X1 U21455 ( .A(n31987), .B(n29324), .C(n14218), .Y(n32269) );
  NAND2X1 U21456 ( .A(n32264), .B(n14371), .Y(n32268) );
  AOI22X1 U21457 ( .A(n32266), .B(n14368), .C(n32265), .D(n14369), .Y(n32267)
         );
  NAND3X1 U21458 ( .A(n32269), .B(n32268), .C(n32267), .Y(n22478) );
  AOI21X1 U21459 ( .A(n30954), .B(n29324), .C(n14218), .Y(n32274) );
  NAND2X1 U21460 ( .A(n32270), .B(n14371), .Y(n32273) );
  AOI22X1 U21461 ( .A(n23325), .B(n14368), .C(n32271), .D(n14369), .Y(n32272)
         );
  NAND3X1 U21462 ( .A(n32274), .B(n32273), .C(n32272), .Y(n22481) );
  AOI21X1 U21463 ( .A(n30975), .B(n29324), .C(n14218), .Y(n32278) );
  NAND2X1 U21464 ( .A(n32275), .B(n14371), .Y(n32277) );
  AOI22X1 U21465 ( .A(n23328), .B(n14368), .C(n23327), .D(n14369), .Y(n32276)
         );
  NAND3X1 U21466 ( .A(n32278), .B(n32277), .C(n32276), .Y(n22484) );
  AOI21X1 U21467 ( .A(n31001), .B(n29324), .C(n14218), .Y(n32282) );
  NAND2X1 U21468 ( .A(n23329), .B(n14371), .Y(n32281) );
  AOI22X1 U21469 ( .A(n23330), .B(n14368), .C(n32279), .D(n14369), .Y(n32280)
         );
  NAND3X1 U21470 ( .A(n32282), .B(n32281), .C(n32280), .Y(n22487) );
  AOI21X1 U21471 ( .A(n31011), .B(n29324), .C(n14218), .Y(n32286) );
  NAND2X1 U21472 ( .A(n32283), .B(n14371), .Y(n32285) );
  AOI22X1 U21473 ( .A(n23333), .B(n14368), .C(n23332), .D(n14369), .Y(n32284)
         );
  NAND3X1 U21474 ( .A(n32286), .B(n32285), .C(n32284), .Y(n22490) );
  AOI21X1 U21475 ( .A(n31038), .B(n29324), .C(n14218), .Y(n32290) );
  NAND2X1 U21476 ( .A(n23334), .B(n14371), .Y(n32289) );
  AOI22X1 U21477 ( .A(n23335), .B(n14368), .C(n32287), .D(n14369), .Y(n32288)
         );
  NAND3X1 U21478 ( .A(n32290), .B(n32289), .C(n32288), .Y(n22493) );
  AOI21X1 U21479 ( .A(n31049), .B(n29324), .C(n14218), .Y(n32294) );
  NAND2X1 U21480 ( .A(n32291), .B(n14371), .Y(n32293) );
  AOI22X1 U21481 ( .A(n23337), .B(n14368), .C(n23336), .D(n14369), .Y(n32292)
         );
  NAND3X1 U21482 ( .A(n32294), .B(n32293), .C(n32292), .Y(n22496) );
  AOI21X1 U21483 ( .A(n31076), .B(n29324), .C(n14218), .Y(n32298) );
  NAND2X1 U21484 ( .A(n23338), .B(n14371), .Y(n32297) );
  AOI22X1 U21485 ( .A(n23339), .B(n14368), .C(n32295), .D(n14369), .Y(n32296)
         );
  NAND3X1 U21486 ( .A(n32298), .B(n32297), .C(n32296), .Y(n22499) );
  AOI21X1 U21487 ( .A(n31089), .B(n29324), .C(n14218), .Y(n32302) );
  NAND2X1 U21488 ( .A(n32299), .B(n14371), .Y(n32301) );
  AOI22X1 U21489 ( .A(n23341), .B(n14368), .C(n23340), .D(n14369), .Y(n32300)
         );
  NAND3X1 U21490 ( .A(n32302), .B(n32301), .C(n32300), .Y(n22502) );
  AOI21X1 U21491 ( .A(n31116), .B(n29324), .C(n14218), .Y(n32306) );
  NAND2X1 U21492 ( .A(n23342), .B(n14371), .Y(n32305) );
  AOI22X1 U21493 ( .A(n23343), .B(n14368), .C(n32303), .D(n14369), .Y(n32304)
         );
  NAND3X1 U21494 ( .A(n32306), .B(n32305), .C(n32304), .Y(n22505) );
  AOI21X1 U21495 ( .A(n31129), .B(n29324), .C(n14218), .Y(n32310) );
  NAND2X1 U21496 ( .A(n32307), .B(n14371), .Y(n32309) );
  AOI22X1 U21497 ( .A(n23345), .B(n14368), .C(n23344), .D(n14369), .Y(n32308)
         );
  NAND3X1 U21498 ( .A(n32310), .B(n32309), .C(n32308), .Y(n22508) );
  AOI21X1 U21499 ( .A(n31156), .B(n29324), .C(n14218), .Y(n32314) );
  NAND2X1 U21500 ( .A(n23346), .B(n14371), .Y(n32313) );
  AOI22X1 U21501 ( .A(n23456), .B(n14368), .C(n32311), .D(n14369), .Y(n32312)
         );
  NAND3X1 U21502 ( .A(n32314), .B(n32313), .C(n32312), .Y(n22511) );
  AOI21X1 U21503 ( .A(n31167), .B(n29325), .C(n14218), .Y(n32318) );
  NAND2X1 U21504 ( .A(n32315), .B(n14371), .Y(n32317) );
  AOI22X1 U21505 ( .A(n23348), .B(n14368), .C(n23347), .D(n14369), .Y(n32316)
         );
  NAND3X1 U21506 ( .A(n32318), .B(n32317), .C(n32316), .Y(n22514) );
  AOI21X1 U21507 ( .A(n31193), .B(n29325), .C(n14218), .Y(n32322) );
  NAND2X1 U21508 ( .A(n23349), .B(n14371), .Y(n32321) );
  AOI22X1 U21509 ( .A(n23350), .B(n14368), .C(n32319), .D(n14369), .Y(n32320)
         );
  NAND3X1 U21510 ( .A(n32322), .B(n32321), .C(n32320), .Y(n22517) );
  AOI21X1 U21511 ( .A(n31206), .B(n29325), .C(n14218), .Y(n32326) );
  NAND2X1 U21512 ( .A(n32323), .B(n14371), .Y(n32325) );
  AOI22X1 U21513 ( .A(n23352), .B(n14368), .C(n23351), .D(n14369), .Y(n32324)
         );
  NAND3X1 U21514 ( .A(n32326), .B(n32325), .C(n32324), .Y(n22520) );
  AOI21X1 U21515 ( .A(n31233), .B(n29325), .C(n14218), .Y(n32330) );
  NAND2X1 U21516 ( .A(n23353), .B(n14371), .Y(n32329) );
  AOI22X1 U21517 ( .A(n23354), .B(n14368), .C(n32327), .D(n14369), .Y(n32328)
         );
  NAND3X1 U21518 ( .A(n32330), .B(n32329), .C(n32328), .Y(n22523) );
  AOI21X1 U21519 ( .A(n31246), .B(n29325), .C(n14218), .Y(n32334) );
  NAND2X1 U21520 ( .A(n32331), .B(n14371), .Y(n32333) );
  AOI22X1 U21521 ( .A(n23356), .B(n14368), .C(n23355), .D(n14369), .Y(n32332)
         );
  NAND3X1 U21522 ( .A(n32334), .B(n32333), .C(n32332), .Y(n22526) );
  AOI21X1 U21523 ( .A(n31273), .B(n29325), .C(n14218), .Y(n32338) );
  NAND2X1 U21524 ( .A(n26274), .B(n14371), .Y(n32337) );
  AOI22X1 U21525 ( .A(n23357), .B(n14368), .C(n32335), .D(n14369), .Y(n32336)
         );
  NAND3X1 U21526 ( .A(n32338), .B(n32337), .C(n32336), .Y(n22529) );
  AOI21X1 U21527 ( .A(n32045), .B(n29325), .C(n14218), .Y(n32342) );
  NAND2X1 U21528 ( .A(n32339), .B(n14371), .Y(n32341) );
  AOI22X1 U21529 ( .A(n23359), .B(n14368), .C(n23358), .D(n14369), .Y(n32340)
         );
  NAND3X1 U21530 ( .A(n32342), .B(n32341), .C(n32340), .Y(n22532) );
  AOI21X1 U21531 ( .A(n31303), .B(n29325), .C(n14218), .Y(n32346) );
  NAND2X1 U21532 ( .A(n32343), .B(n14371), .Y(n32345) );
  AOI22X1 U21533 ( .A(n23361), .B(n14368), .C(n23360), .D(n14369), .Y(n32344)
         );
  NAND3X1 U21534 ( .A(n32346), .B(n32345), .C(n32344), .Y(n22535) );
  AOI21X1 U21535 ( .A(n32053), .B(n29325), .C(n14218), .Y(n32350) );
  NAND2X1 U21536 ( .A(n32347), .B(n14371), .Y(n32349) );
  AOI22X1 U21537 ( .A(n23363), .B(n14368), .C(n23362), .D(n14369), .Y(n32348)
         );
  NAND3X1 U21538 ( .A(n32350), .B(n32349), .C(n32348), .Y(n22538) );
  AOI21X1 U21539 ( .A(n31340), .B(n29325), .C(n14218), .Y(n32354) );
  NAND2X1 U21540 ( .A(n32351), .B(n14371), .Y(n32353) );
  AOI22X1 U21541 ( .A(n23366), .B(n14368), .C(n23365), .D(n14369), .Y(n32352)
         );
  NAND3X1 U21542 ( .A(n32354), .B(n32353), .C(n32352), .Y(n22541) );
  AOI21X1 U21543 ( .A(n32060), .B(n29325), .C(n14218), .Y(n32358) );
  NAND2X1 U21544 ( .A(n32355), .B(n14371), .Y(n32357) );
  AOI22X1 U21545 ( .A(n23368), .B(n14368), .C(n23367), .D(n14369), .Y(n32356)
         );
  NAND3X1 U21546 ( .A(n32358), .B(n32357), .C(n32356), .Y(n22544) );
  AOI21X1 U21547 ( .A(n31380), .B(n29325), .C(n14218), .Y(n32362) );
  NAND2X1 U21548 ( .A(n32359), .B(n14371), .Y(n32361) );
  AOI22X1 U21549 ( .A(n23370), .B(n14368), .C(n23369), .D(n14369), .Y(n32360)
         );
  NAND3X1 U21550 ( .A(n32362), .B(n32361), .C(n32360), .Y(n22547) );
  AOI21X1 U21551 ( .A(n32068), .B(n29325), .C(n14218), .Y(n32366) );
  NAND2X1 U21552 ( .A(n32363), .B(n14371), .Y(n32365) );
  AOI22X1 U21553 ( .A(n23372), .B(n14368), .C(n23371), .D(n14369), .Y(n32364)
         );
  NAND3X1 U21554 ( .A(n32366), .B(n32365), .C(n32364), .Y(n22550) );
  AOI21X1 U21555 ( .A(n31421), .B(n29326), .C(n14218), .Y(n32370) );
  NAND2X1 U21556 ( .A(n32367), .B(n14371), .Y(n32369) );
  AOI22X1 U21557 ( .A(n23374), .B(n14368), .C(n23373), .D(n14369), .Y(n32368)
         );
  NAND3X1 U21558 ( .A(n32370), .B(n32369), .C(n32368), .Y(n22553) );
  AOI21X1 U21559 ( .A(n32076), .B(n29326), .C(n14218), .Y(n32374) );
  NAND2X1 U21560 ( .A(n32371), .B(n14371), .Y(n32373) );
  AOI22X1 U21561 ( .A(n23376), .B(n14368), .C(n23375), .D(n14369), .Y(n32372)
         );
  NAND3X1 U21562 ( .A(n32374), .B(n32373), .C(n32372), .Y(n22556) );
  AOI21X1 U21563 ( .A(n31460), .B(n29326), .C(n14218), .Y(n32378) );
  NAND2X1 U21564 ( .A(n32375), .B(n14371), .Y(n32377) );
  AOI22X1 U21565 ( .A(n23378), .B(n14368), .C(n23377), .D(n14369), .Y(n32376)
         );
  NAND3X1 U21566 ( .A(n32378), .B(n32377), .C(n32376), .Y(n22559) );
  AOI21X1 U21567 ( .A(n32084), .B(n29326), .C(n14218), .Y(n32382) );
  NAND2X1 U21568 ( .A(n32379), .B(n14371), .Y(n32381) );
  AOI22X1 U21569 ( .A(n23380), .B(n14368), .C(n23379), .D(n14369), .Y(n32380)
         );
  NAND3X1 U21570 ( .A(n32382), .B(n32381), .C(n32380), .Y(n22562) );
  AOI21X1 U21571 ( .A(n31499), .B(n29326), .C(n14218), .Y(n32386) );
  NAND2X1 U21572 ( .A(n32383), .B(n14371), .Y(n32385) );
  AOI22X1 U21573 ( .A(n23383), .B(n14368), .C(n23382), .D(n14369), .Y(n32384)
         );
  NAND3X1 U21574 ( .A(n32386), .B(n32385), .C(n32384), .Y(n22565) );
  AOI21X1 U21575 ( .A(n32091), .B(n29326), .C(n14218), .Y(n32390) );
  NAND2X1 U21576 ( .A(n32387), .B(n14371), .Y(n32389) );
  AOI22X1 U21577 ( .A(n23385), .B(n14368), .C(n23384), .D(n14369), .Y(n32388)
         );
  NAND3X1 U21578 ( .A(n32390), .B(n32389), .C(n32388), .Y(n22568) );
  AOI21X1 U21579 ( .A(n31537), .B(n29326), .C(n14218), .Y(n32394) );
  NAND2X1 U21580 ( .A(n32391), .B(n14371), .Y(n32393) );
  AOI22X1 U21581 ( .A(n23387), .B(n14368), .C(n23386), .D(n14369), .Y(n32392)
         );
  NAND3X1 U21582 ( .A(n32394), .B(n32393), .C(n32392), .Y(n22571) );
  AOI21X1 U21583 ( .A(n32100), .B(n29326), .C(n14218), .Y(n32398) );
  NAND2X1 U21584 ( .A(n32395), .B(n14371), .Y(n32397) );
  AOI22X1 U21585 ( .A(n23389), .B(n14368), .C(n23388), .D(n14369), .Y(n32396)
         );
  NAND3X1 U21586 ( .A(n32398), .B(n32397), .C(n32396), .Y(n22574) );
  AOI21X1 U21587 ( .A(n31578), .B(n29326), .C(n14218), .Y(n32402) );
  NAND2X1 U21588 ( .A(n32399), .B(n14371), .Y(n32401) );
  AOI22X1 U21589 ( .A(n23391), .B(n14368), .C(n23390), .D(n14369), .Y(n32400)
         );
  NAND3X1 U21590 ( .A(n32402), .B(n32401), .C(n32400), .Y(n22577) );
  AOI21X1 U21591 ( .A(n31598), .B(n29326), .C(n14218), .Y(n32406) );
  NAND2X1 U21592 ( .A(n32403), .B(n14371), .Y(n32405) );
  AOI22X1 U21593 ( .A(n23393), .B(n14368), .C(n23392), .D(n14369), .Y(n32404)
         );
  NAND3X1 U21594 ( .A(n32406), .B(n32405), .C(n32404), .Y(n22580) );
  AOI21X1 U21595 ( .A(n31624), .B(n29326), .C(n14218), .Y(n32410) );
  NAND2X1 U21596 ( .A(n23394), .B(n14371), .Y(n32409) );
  AOI22X1 U21597 ( .A(n23395), .B(n14368), .C(n32407), .D(n14369), .Y(n32408)
         );
  NAND3X1 U21598 ( .A(n32410), .B(n32409), .C(n32408), .Y(n22583) );
  AOI21X1 U21599 ( .A(n31635), .B(n29326), .C(n14218), .Y(n32414) );
  NAND2X1 U21600 ( .A(n32411), .B(n14371), .Y(n32413) );
  AOI22X1 U21601 ( .A(n23397), .B(n14368), .C(n23396), .D(n14369), .Y(n32412)
         );
  NAND3X1 U21602 ( .A(n32414), .B(n32413), .C(n32412), .Y(n22586) );
  AOI21X1 U21603 ( .A(n31660), .B(n29326), .C(n14218), .Y(n32418) );
  NAND2X1 U21604 ( .A(n23398), .B(n14371), .Y(n32417) );
  AOI22X1 U21605 ( .A(n23399), .B(n14368), .C(n32415), .D(n14369), .Y(n32416)
         );
  NAND3X1 U21606 ( .A(n32418), .B(n32417), .C(n32416), .Y(n22589) );
  AOI21X1 U21607 ( .A(n31672), .B(n29327), .C(n14218), .Y(n32422) );
  NAND2X1 U21608 ( .A(n32419), .B(n14371), .Y(n32421) );
  AOI22X1 U21609 ( .A(n23401), .B(n14368), .C(n23400), .D(n14369), .Y(n32420)
         );
  NAND3X1 U21610 ( .A(n32422), .B(n32421), .C(n32420), .Y(n22592) );
  AOI21X1 U21611 ( .A(n31698), .B(n29327), .C(n14218), .Y(n32426) );
  NAND2X1 U21612 ( .A(n23402), .B(n14371), .Y(n32425) );
  AOI22X1 U21613 ( .A(n23403), .B(n14368), .C(n32423), .D(n14369), .Y(n32424)
         );
  NAND3X1 U21614 ( .A(n32426), .B(n32425), .C(n32424), .Y(n22595) );
  AOI21X1 U21615 ( .A(n31711), .B(n29327), .C(n14218), .Y(n32430) );
  NAND2X1 U21616 ( .A(n32427), .B(n14371), .Y(n32429) );
  AOI22X1 U21617 ( .A(n23405), .B(n14368), .C(n23404), .D(n14369), .Y(n32428)
         );
  NAND3X1 U21618 ( .A(n32430), .B(n32429), .C(n32428), .Y(n22598) );
  AOI21X1 U21619 ( .A(n31738), .B(n29327), .C(n14218), .Y(n32433) );
  NAND2X1 U21620 ( .A(n23406), .B(n14371), .Y(n32432) );
  AOI22X1 U21621 ( .A(n23408), .B(n14368), .C(n23407), .D(n14369), .Y(n32431)
         );
  NAND3X1 U21622 ( .A(n32433), .B(n32432), .C(n32431), .Y(n22601) );
  AOI21X1 U21623 ( .A(n31749), .B(n29327), .C(n14218), .Y(n32437) );
  NAND2X1 U21624 ( .A(n32434), .B(n14371), .Y(n32436) );
  AOI22X1 U21625 ( .A(n23410), .B(n14368), .C(n23409), .D(n14369), .Y(n32435)
         );
  NAND3X1 U21626 ( .A(n32437), .B(n32436), .C(n32435), .Y(n22604) );
  AOI21X1 U21627 ( .A(n31776), .B(n29327), .C(n14218), .Y(n32441) );
  NAND2X1 U21628 ( .A(n23411), .B(n14371), .Y(n32440) );
  AOI22X1 U21629 ( .A(n23412), .B(n14368), .C(n32438), .D(n14369), .Y(n32439)
         );
  NAND3X1 U21630 ( .A(n32441), .B(n32440), .C(n32439), .Y(n22607) );
  AOI21X1 U21631 ( .A(n31789), .B(n29327), .C(n14218), .Y(n32445) );
  NAND2X1 U21632 ( .A(n32442), .B(n14371), .Y(n32444) );
  AOI22X1 U21633 ( .A(n23414), .B(n14368), .C(n23413), .D(n14369), .Y(n32443)
         );
  NAND3X1 U21634 ( .A(n32445), .B(n32444), .C(n32443), .Y(n22610) );
  AOI21X1 U21635 ( .A(n31815), .B(n29327), .C(n14218), .Y(n32449) );
  NAND2X1 U21636 ( .A(n23415), .B(n14371), .Y(n32448) );
  AOI22X1 U21637 ( .A(n23416), .B(n14368), .C(n32446), .D(n14369), .Y(n32447)
         );
  NAND3X1 U21638 ( .A(n32449), .B(n32448), .C(n32447), .Y(n22613) );
  AOI21X1 U21639 ( .A(n31828), .B(n29327), .C(n14218), .Y(n32453) );
  NAND2X1 U21640 ( .A(n32450), .B(n14371), .Y(n32452) );
  AOI22X1 U21641 ( .A(n23418), .B(n14368), .C(n23417), .D(n14369), .Y(n32451)
         );
  NAND3X1 U21642 ( .A(n32453), .B(n32452), .C(n32451), .Y(n22616) );
  AOI21X1 U21643 ( .A(n31855), .B(n29327), .C(n14218), .Y(n32456) );
  NAND2X1 U21644 ( .A(n23419), .B(n14371), .Y(n32455) );
  AOI22X1 U21645 ( .A(n23421), .B(n14368), .C(n23420), .D(n14369), .Y(n32454)
         );
  NAND3X1 U21646 ( .A(n32456), .B(n32455), .C(n32454), .Y(n22619) );
  AOI21X1 U21647 ( .A(n31867), .B(n29327), .C(n14218), .Y(n32460) );
  NAND2X1 U21648 ( .A(n32457), .B(n14371), .Y(n32459) );
  AOI22X1 U21649 ( .A(n14368), .B(n23423), .C(n14369), .D(n23422), .Y(n32458)
         );
  NAND3X1 U21650 ( .A(n32460), .B(n32459), .C(n32458), .Y(n22622) );
  NAND2X1 U21651 ( .A(n29327), .B(n32461), .Y(n32465) );
  AOI21X1 U21652 ( .A(n14371), .B(n32463), .C(n14218), .Y(n32464) );
  NAND3X1 U21653 ( .A(n14366), .B(n32465), .C(n32464), .Y(n22625) );
  AOI22X1 U21654 ( .A(n3154), .B(n29836), .C(n3148), .D(n29824), .Y(n32466) );
  OAI21X1 U21655 ( .A(n27206), .B(n32696), .C(n21573), .Y(n32470) );
  AOI22X1 U21656 ( .A(n3136), .B(n25769), .C(n3130), .D(n29794), .Y(n32467) );
  OAI21X1 U21657 ( .A(n27025), .B(n32468), .C(n21574), .Y(n32469) );
  AOI22X1 U21658 ( .A(n3166), .B(n26519), .C(n3160), .D(n23450), .Y(n32471) );
  OAI21X1 U21659 ( .A(n27119), .B(n32472), .C(n21575), .Y(n32476) );
  AOI22X1 U21660 ( .A(n3184), .B(n33019), .C(n3178), .D(n26518), .Y(n32473) );
  OAI21X1 U21661 ( .A(n27024), .B(n32474), .C(n21576), .Y(n32475) );
  AOI22X1 U21662 ( .A(n3242), .B(n32477), .C(n3254), .D(n32478), .Y(n32483) );
  AOI22X1 U21663 ( .A(n3266), .B(n23455), .C(n3224), .D(n32480), .Y(n32481) );
  NAND3X1 U21664 ( .A(n22500), .B(n21490), .C(n24779), .Y(n32488) );
  AOI22X1 U21665 ( .A(n3118), .B(n25830), .C(n3248), .D(n32957), .Y(n32484) );
  OAI21X1 U21666 ( .A(n25443), .B(n33373), .C(n21577), .Y(n32487) );
  AOI22X1 U21667 ( .A(n3106), .B(n33884), .C(RO[176]), .D(n27250), .Y(n32485)
         );
  OAI21X1 U21668 ( .A(n27189), .B(n33185), .C(n21578), .Y(n32486) );
  NOR3X1 U21669 ( .A(n22882), .B(n32487), .C(n32486), .Y(n32513) );
  AOI22X1 U21670 ( .A(n3176), .B(n27225), .C(n3188), .D(n23470), .Y(n32494) );
  AOI22X1 U21671 ( .A(n32490), .B(n25696), .C(RO[178]), .D(n27298), .Y(n32492)
         );
  NAND3X1 U21672 ( .A(n22503), .B(n21493), .C(n22748), .Y(n32501) );
  AOI22X1 U21673 ( .A(n3230), .B(n25491), .C(n3182), .D(n32783), .Y(n32495) );
  OAI21X1 U21674 ( .A(n27078), .B(n32496), .C(n21579), .Y(n32500) );
  AOI22X1 U21675 ( .A(n3218), .B(n23307), .C(n3212), .D(n23306), .Y(n32497) );
  OAI21X1 U21676 ( .A(n21222), .B(n32498), .C(n21580), .Y(n32499) );
  NOR3X1 U21677 ( .A(n32499), .B(n32500), .C(n24919), .Y(n32511) );
  AOI22X1 U21678 ( .A(n3134), .B(n32988), .C(n3140), .D(n21139), .Y(n32504) );
  AOI22X1 U21679 ( .A(n3158), .B(n27232), .C(n3164), .D(n21220), .Y(n32502) );
  AOI22X1 U21680 ( .A(n3122), .B(n27219), .C(n3104), .D(n27217), .Y(n32505) );
  OAI21X1 U21681 ( .A(n26996), .B(n32506), .C(n21581), .Y(n32509) );
  AOI22X1 U21682 ( .A(n3128), .B(n27220), .C(n3116), .D(n27216), .Y(n32507) );
  OAI21X1 U21683 ( .A(n27115), .B(n32567), .C(n21582), .Y(n32508) );
  NOR3X1 U21684 ( .A(n32508), .B(n32509), .C(n22883), .Y(n32510) );
  NAND3X1 U21685 ( .A(n32514), .B(n32513), .C(n32512), .Y(n32515) );
  AOI22X1 U21686 ( .A(n3108), .B(n33875), .C(n33900), .D(n3102), .Y(n32516) );
  OAI21X1 U21687 ( .A(n26269), .B(n32517), .C(n21583), .Y(n32521) );
  AOI22X1 U21688 ( .A(n3268), .B(n33216), .C(n3262), .D(n33247), .Y(n32519) );
  OAI21X1 U21689 ( .A(n21375), .B(n32659), .C(n21584), .Y(n32520) );
  AOI22X1 U21690 ( .A(n3126), .B(n33806), .C(n25675), .D(n3120), .Y(n32522) );
  OAI21X1 U21691 ( .A(n27199), .B(n32523), .C(n21585), .Y(n32526) );
  AOI22X1 U21692 ( .A(n3144), .B(n26077), .C(n3138), .D(n33762), .Y(n32524) );
  OAI21X1 U21693 ( .A(n21378), .B(n32602), .C(n21586), .Y(n32525) );
  NOR3X1 U21694 ( .A(n32527), .B(n32526), .C(n32525), .Y(n32564) );
  AOI22X1 U21695 ( .A(n3196), .B(n33538), .C(n3190), .D(n33560), .Y(n32532) );
  AOI22X1 U21696 ( .A(n3220), .B(n33912), .C(n3214), .D(n33471), .Y(n32530) );
  NAND3X1 U21697 ( .A(n22506), .B(n21496), .C(n24781), .Y(n32540) );
  AOI22X1 U21698 ( .A(n3232), .B(n33399), .C(n3226), .D(n33430), .Y(n32534) );
  OAI21X1 U21699 ( .A(n25452), .B(n32535), .C(n21587), .Y(n32539) );
  AOI22X1 U21700 ( .A(n3250), .B(n33308), .C(n3244), .D(n33339), .Y(n32537) );
  OAI21X1 U21701 ( .A(n25454), .B(n32687), .C(n21588), .Y(n32538) );
  NOR3X1 U21702 ( .A(n22887), .B(n32539), .C(n32538), .Y(n32563) );
  AOI22X1 U21703 ( .A(n3222), .B(n33429), .C(n3216), .D(n33462), .Y(n32543) );
  AOI22X1 U21704 ( .A(n3240), .B(n25680), .C(n3234), .D(n25657), .Y(n32541) );
  AOI22X1 U21705 ( .A(n3258), .B(n25658), .C(n3252), .D(n33295), .Y(n32544) );
  OAI21X1 U21706 ( .A(n21384), .B(n32582), .C(n21589), .Y(n32548) );
  AOI22X1 U21707 ( .A(RO[174]), .B(n23457), .C(n3270), .D(n34222), .Y(n32545)
         );
  OAI21X1 U21708 ( .A(n21387), .B(n32546), .C(n21590), .Y(n32547) );
  NOR3X1 U21709 ( .A(n22928), .B(n32548), .C(n32547), .Y(n32561) );
  AOI22X1 U21710 ( .A(n3156), .B(n33696), .C(n3150), .D(n33718), .Y(n32552) );
  AOI22X1 U21711 ( .A(n3174), .B(n21232), .C(n3168), .D(n33653), .Y(n32550) );
  NAND3X1 U21712 ( .A(n24123), .B(n24589), .C(n22749), .Y(n32559) );
  AOI22X1 U21713 ( .A(n3192), .B(n33551), .C(n3186), .D(n33587), .Y(n32554) );
  OAI21X1 U21714 ( .A(n27207), .B(n32593), .C(n21591), .Y(n32558) );
  AOI22X1 U21715 ( .A(n3210), .B(n33485), .C(n3204), .D(n33508), .Y(n32555) );
  OAI21X1 U21716 ( .A(n25457), .B(n32556), .C(n21592), .Y(n32557) );
  NOR3X1 U21717 ( .A(n22888), .B(n32558), .C(n32557), .Y(n32560) );
  NAND3X1 U21718 ( .A(n32564), .B(n32563), .C(n32562), .Y(n32565) );
  AOI22X1 U21719 ( .A(n3146), .B(n29824), .C(n3134), .D(n25769), .Y(n32566) );
  OAI21X1 U21720 ( .A(n27204), .B(n32567), .C(n21593), .Y(n32571) );
  AOI22X1 U21721 ( .A(n3116), .B(n29190), .C(n3128), .D(n29794), .Y(n32568) );
  OAI21X1 U21722 ( .A(n27026), .B(n32569), .C(n21594), .Y(n32570) );
  AOI22X1 U21723 ( .A(n23450), .B(n3158), .C(n3152), .D(n29836), .Y(n32572) );
  OAI21X1 U21724 ( .A(n27121), .B(n32573), .C(n21595), .Y(n32576) );
  AOI22X1 U21725 ( .A(n3176), .B(n26518), .C(n3170), .D(n33639), .Y(n32574) );
  OAI21X1 U21726 ( .A(n32953), .B(n32740), .C(n21596), .Y(n32575) );
  NOR3X1 U21727 ( .A(n32576), .B(n32575), .C(n32577), .Y(n32611) );
  AOI22X1 U21728 ( .A(n3240), .B(n32477), .C(n3252), .D(n32478), .Y(n32580) );
  AOI22X1 U21729 ( .A(n3258), .B(n23451), .C(n3222), .D(n32480), .Y(n32578) );
  AOI22X1 U21730 ( .A(n3264), .B(n23453), .C(n3234), .D(n32961), .Y(n32581) );
  OAI21X1 U21731 ( .A(n32964), .B(n32582), .C(n21597), .Y(n32586) );
  AOI22X1 U21732 ( .A(n3104), .B(n33884), .C(RO[174]), .D(n27250), .Y(n32583)
         );
  OAI21X1 U21733 ( .A(n27189), .B(n32584), .C(n21598), .Y(n32585) );
  NOR3X1 U21734 ( .A(n32585), .B(n32586), .C(n22889), .Y(n32610) );
  AOI22X1 U21735 ( .A(n3174), .B(n27225), .C(n3186), .D(n23470), .Y(n32591) );
  AOI22X1 U21736 ( .A(n3192), .B(n23471), .C(n27048), .D(n29933), .Y(n32589)
         );
  AOI22X1 U21737 ( .A(n3198), .B(n32490), .C(n3168), .D(n32871), .Y(n32592) );
  OAI21X1 U21738 ( .A(n26870), .B(n32593), .C(n21666), .Y(n32596) );
  AOI22X1 U21739 ( .A(n3216), .B(n23307), .C(n3210), .D(n23306), .Y(n32594) );
  OAI21X1 U21740 ( .A(n21222), .B(n32722), .C(n21699), .Y(n32595) );
  NOR3X1 U21741 ( .A(n32596), .B(n32597), .C(n32595), .Y(n32608) );
  AOI22X1 U21742 ( .A(n3126), .B(n27220), .C(n3138), .D(n27218), .Y(n32600) );
  AOI22X1 U21743 ( .A(n3144), .B(n32882), .C(n3156), .D(n27232), .Y(n32598) );
  AOI22X1 U21744 ( .A(n3120), .B(n27219), .C(n3102), .D(n27217), .Y(n32601) );
  OAI21X1 U21745 ( .A(n26931), .B(n32602), .C(n21767), .Y(n32606) );
  AOI22X1 U21746 ( .A(RO[176]), .B(n27298), .C(n3114), .D(n27216), .Y(n32603)
         );
  OAI21X1 U21747 ( .A(n27115), .B(n32604), .C(n21782), .Y(n32605) );
  NOR3X1 U21748 ( .A(n22893), .B(n32606), .C(n32605), .Y(n32607) );
  NAND3X1 U21749 ( .A(n32610), .B(n32611), .C(n32609), .Y(n32612) );
  AOI22X1 U21750 ( .A(n33852), .B(n3112), .C(n3106), .D(n33875), .Y(n32613) );
  OAI21X1 U21751 ( .A(n25442), .B(n33312), .C(n21801), .Y(n32616) );
  AOI22X1 U21752 ( .A(n3260), .B(n33247), .C(n3254), .D(n33277), .Y(n32614) );
  OAI21X1 U21753 ( .A(n27200), .B(n33185), .C(n21848), .Y(n32615) );
  AOI22X1 U21754 ( .A(n3124), .B(n33806), .C(n3118), .D(n25675), .Y(n32617) );
  OAI21X1 U21755 ( .A(n27195), .B(n33220), .C(n21849), .Y(n32621) );
  AOI22X1 U21756 ( .A(n3142), .B(n26077), .C(n3136), .D(n33762), .Y(n32618) );
  OAI21X1 U21757 ( .A(n21378), .B(n32619), .C(n21850), .Y(n32620) );
  NOR3X1 U21758 ( .A(n32620), .B(n32621), .C(n32622), .Y(n32656) );
  AOI22X1 U21759 ( .A(n3194), .B(n33538), .C(n3188), .D(n33560), .Y(n32625) );
  AOI22X1 U21760 ( .A(n3212), .B(n33471), .C(n33517), .D(n25775), .Y(n32623)
         );
  NAND3X1 U21761 ( .A(n22509), .B(n24590), .C(n24783), .Y(n32631) );
  AOI22X1 U21762 ( .A(n3224), .B(n33430), .C(n3218), .D(n33912), .Y(n32626) );
  OAI21X1 U21763 ( .A(n26078), .B(n32627), .C(n21851), .Y(n32630) );
  AOI22X1 U21764 ( .A(n3242), .B(n33339), .C(n3236), .D(n33369), .Y(n32628) );
  OAI21X1 U21765 ( .A(n21435), .B(n33403), .C(n23774), .Y(n32629) );
  NOR3X1 U21766 ( .A(n32629), .B(n32630), .C(n23616), .Y(n32655) );
  AOI22X1 U21767 ( .A(n3220), .B(n33429), .C(n3214), .D(n33462), .Y(n32634) );
  AOI22X1 U21768 ( .A(n3238), .B(n25680), .C(n3232), .D(n25657), .Y(n32632) );
  AOI22X1 U21769 ( .A(n3256), .B(n25658), .C(n3250), .D(n33295), .Y(n32635) );
  OAI21X1 U21770 ( .A(n21384), .B(n32636), .C(n23775), .Y(n32640) );
  AOI22X1 U21771 ( .A(n3274), .B(n23457), .C(n3268), .D(n34222), .Y(n32637) );
  OAI21X1 U21772 ( .A(n21387), .B(n32638), .C(n21853), .Y(n32639) );
  NOR3X1 U21773 ( .A(n32639), .B(n32640), .C(n22929), .Y(n32653) );
  AOI22X1 U21774 ( .A(n33696), .B(n3154), .C(n3148), .D(n33718), .Y(n32644) );
  AOI22X1 U21775 ( .A(n3172), .B(n21232), .C(n3166), .D(n33653), .Y(n32642) );
  NAND3X1 U21776 ( .A(n22512), .B(n21499), .C(n24785), .Y(n32651) );
  AOI22X1 U21777 ( .A(n3190), .B(n33551), .C(n3184), .D(n33587), .Y(n32645) );
  OAI21X1 U21778 ( .A(n27207), .B(n32646), .C(n21855), .Y(n32650) );
  AOI22X1 U21779 ( .A(n3208), .B(n33485), .C(n3202), .D(n33508), .Y(n32647) );
  OAI21X1 U21780 ( .A(n25456), .B(n32648), .C(n21856), .Y(n32649) );
  NOR3X1 U21781 ( .A(n32649), .B(n32650), .C(n24921), .Y(n32652) );
  NAND3X1 U21782 ( .A(n32656), .B(n32654), .C(n32655), .Y(n32657) );
  AOI22X1 U21783 ( .A(n3156), .B(n29836), .C(n3150), .D(n29824), .Y(n32658) );
  OAI21X1 U21784 ( .A(n27204), .B(n32659), .C(n21857), .Y(n32663) );
  AOI22X1 U21785 ( .A(n3138), .B(n29803), .C(n3132), .D(n29794), .Y(n32660) );
  OAI21X1 U21786 ( .A(n27027), .B(n32661), .C(n21859), .Y(n32662) );
  AOI22X1 U21787 ( .A(n3168), .B(n26519), .C(n3162), .D(n23450), .Y(n32664) );
  OAI21X1 U21788 ( .A(n27121), .B(n32665), .C(n21861), .Y(n32669) );
  AOI22X1 U21789 ( .A(n3186), .B(n26520), .C(n3180), .D(n26518), .Y(n32666) );
  OAI21X1 U21790 ( .A(n27024), .B(n32667), .C(n21862), .Y(n32668) );
  NOR3X1 U21791 ( .A(n32670), .B(n32669), .C(n32668), .Y(n32703) );
  AOI22X1 U21792 ( .A(n3244), .B(n32477), .C(n3262), .D(n23451), .Y(n32673) );
  AOI22X1 U21793 ( .A(n3268), .B(n23455), .C(n3226), .D(n32480), .Y(n32671) );
  NAND3X1 U21794 ( .A(n24787), .B(n21502), .C(n22515), .Y(n32680) );
  AOI22X1 U21795 ( .A(n33908), .B(n3102), .C(n3256), .D(n32478), .Y(n32674) );
  OAI21X1 U21796 ( .A(n25394), .B(n32675), .C(n21863), .Y(n32679) );
  AOI22X1 U21797 ( .A(n3108), .B(n33884), .C(RO[178]), .D(n27250), .Y(n32676)
         );
  OAI21X1 U21798 ( .A(n32773), .B(n32677), .C(n21864), .Y(n32678) );
  NOR3X1 U21799 ( .A(n32678), .B(n32679), .C(n22896), .Y(n32702) );
  AOI22X1 U21800 ( .A(n3178), .B(n27225), .C(n3196), .D(n23471), .Y(n32683) );
  AOI22X1 U21801 ( .A(n3202), .B(n32490), .C(n3136), .D(n32988), .Y(n32681) );
  AOI22X1 U21802 ( .A(n3232), .B(n25491), .C(n3190), .D(n23470), .Y(n32684) );
  OAI21X1 U21803 ( .A(n25404), .B(n32685), .C(n21865), .Y(n32689) );
  AOI22X1 U21804 ( .A(n3220), .B(n23307), .C(n3214), .D(n23306), .Y(n32686) );
  OAI21X1 U21805 ( .A(n25444), .B(n32687), .C(n21866), .Y(n32688) );
  NOR3X1 U21806 ( .A(n22897), .B(n32689), .C(n32688), .Y(n32700) );
  AOI22X1 U21807 ( .A(n3148), .B(n21188), .C(n3142), .D(n27218), .Y(n32692) );
  AOI22X1 U21808 ( .A(n3172), .B(n21152), .C(n3166), .D(n32877), .Y(n32690) );
  AOI22X1 U21809 ( .A(n27219), .B(n3124), .C(n3106), .D(n27217), .Y(n32693) );
  OAI21X1 U21810 ( .A(n32694), .B(n26811), .C(n21867), .Y(n32698) );
  AOI22X1 U21811 ( .A(n3130), .B(n27220), .C(n3118), .D(n27216), .Y(n32695) );
  OAI21X1 U21812 ( .A(n27115), .B(n32696), .C(n21868), .Y(n32697) );
  NOR3X1 U21813 ( .A(n22901), .B(n32697), .C(n32698), .Y(n32699) );
  NAND3X1 U21814 ( .A(n32703), .B(n32702), .C(n32701), .Y(n32704) );
  AOI22X1 U21815 ( .A(n33875), .B(n3110), .C(n33900), .D(n3104), .Y(n32705) );
  OAI21X1 U21816 ( .A(n26269), .B(n32706), .C(n21869), .Y(n32710) );
  OAI21X1 U21817 ( .A(n21375), .B(n32708), .C(n21870), .Y(n32709) );
  AOI22X1 U21818 ( .A(n3128), .B(n33806), .C(n3122), .D(n33829), .Y(n32711) );
  OAI21X1 U21819 ( .A(n27198), .B(n32712), .C(n21871), .Y(n32716) );
  AOI22X1 U21820 ( .A(n3146), .B(n26077), .C(n3140), .D(n33762), .Y(n32713) );
  OAI21X1 U21821 ( .A(n21378), .B(n32714), .C(n23776), .Y(n32715) );
  NOR3X1 U21822 ( .A(n32717), .B(n32716), .C(n32715), .Y(n32750) );
  AOI22X1 U21823 ( .A(n3198), .B(n25628), .C(n3192), .D(n33560), .Y(n32720) );
  AOI22X1 U21824 ( .A(n3222), .B(n33912), .C(n3216), .D(n33471), .Y(n32718) );
  NAND3X1 U21825 ( .A(n22518), .B(n21505), .C(n24789), .Y(n32727) );
  AOI22X1 U21826 ( .A(n3234), .B(n33399), .C(n3228), .D(n33430), .Y(n32721) );
  OAI21X1 U21827 ( .A(n25452), .B(n32722), .C(n21872), .Y(n32726) );
  AOI22X1 U21828 ( .A(n3252), .B(n33308), .C(n3246), .D(n33339), .Y(n32723) );
  OAI21X1 U21829 ( .A(n25454), .B(n32724), .C(n23777), .Y(n32725) );
  NOR3X1 U21830 ( .A(n32725), .B(n32726), .C(n22905), .Y(n32749) );
  AOI22X1 U21831 ( .A(n3224), .B(n33429), .C(n3218), .D(n33462), .Y(n32730) );
  AOI22X1 U21832 ( .A(n3242), .B(n25680), .C(n3236), .D(n25657), .Y(n32728) );
  AOI22X1 U21833 ( .A(n3260), .B(n25658), .C(n3254), .D(n33295), .Y(n32731) );
  OAI21X1 U21834 ( .A(n21384), .B(n33403), .C(n21873), .Y(n32734) );
  AOI22X1 U21835 ( .A(RO[176]), .B(n23457), .C(n3272), .D(n34222), .Y(n32732)
         );
  OAI21X1 U21836 ( .A(n21387), .B(n33220), .C(n21874), .Y(n32733) );
  NOR3X1 U21837 ( .A(n32735), .B(n32734), .C(n32733), .Y(n32747) );
  AOI22X1 U21838 ( .A(n3158), .B(n33696), .C(n3152), .D(n33718), .Y(n32738) );
  AOI22X1 U21839 ( .A(n3176), .B(n21232), .C(n3170), .D(n33653), .Y(n32736) );
  AOI22X1 U21840 ( .A(n3194), .B(n33551), .C(n3188), .D(n33587), .Y(n32739) );
  OAI21X1 U21841 ( .A(n27207), .B(n32740), .C(n21875), .Y(n32744) );
  AOI22X1 U21842 ( .A(n3212), .B(n33485), .C(n3206), .D(n33508), .Y(n32741) );
  OAI21X1 U21843 ( .A(n32742), .B(n25456), .C(n21876), .Y(n32743) );
  NOR3X1 U21844 ( .A(n32744), .B(n32745), .C(n32743), .Y(n32746) );
  AND2X2 U21845 ( .A(n32747), .B(n32746), .Y(n32748) );
  NAND3X1 U21846 ( .A(n32750), .B(n32749), .C(n32748), .Y(n32751) );
  AOI22X1 U21847 ( .A(n3157), .B(n29836), .C(n3151), .D(n29824), .Y(n32752) );
  OAI21X1 U21848 ( .A(n27203), .B(n32897), .C(n21877), .Y(n32756) );
  AOI22X1 U21849 ( .A(n3139), .B(n29803), .C(n3133), .D(n29794), .Y(n32753) );
  OAI21X1 U21850 ( .A(n27025), .B(n32754), .C(n21878), .Y(n32755) );
  AOI22X1 U21851 ( .A(n3169), .B(n26519), .C(n3163), .D(n23450), .Y(n32757) );
  OAI21X1 U21852 ( .A(n27119), .B(n32758), .C(n21879), .Y(n32762) );
  AOI22X1 U21853 ( .A(n33019), .B(n3187), .C(n3181), .D(n26518), .Y(n32759) );
  OAI21X1 U21854 ( .A(n27023), .B(n32760), .C(n21880), .Y(n32761) );
  NOR3X1 U21855 ( .A(n32761), .B(n32762), .C(n32763), .Y(n32800) );
  AOI22X1 U21856 ( .A(n3245), .B(n32477), .C(n3263), .D(n23451), .Y(n32767) );
  AOI22X1 U21857 ( .A(n3269), .B(n23454), .C(n3227), .D(n32480), .Y(n32765) );
  NAND3X1 U21858 ( .A(n22521), .B(n22731), .C(n22750), .Y(n32776) );
  AOI22X1 U21859 ( .A(n33908), .B(n3103), .C(n3257), .D(n32478), .Y(n32768) );
  OAI21X1 U21860 ( .A(n25394), .B(n32769), .C(n21881), .Y(n32775) );
  AOI22X1 U21861 ( .A(n25751), .B(n33884), .C(RO[179]), .D(n27250), .Y(n32771)
         );
  OAI21X1 U21862 ( .A(n32773), .B(n32772), .C(n21882), .Y(n32774) );
  NOR3X1 U21863 ( .A(n24883), .B(n32775), .C(n32774), .Y(n32799) );
  AOI22X1 U21864 ( .A(n3179), .B(n27225), .C(n3197), .D(n32973), .Y(n32780) );
  AOI22X1 U21865 ( .A(n3203), .B(n32490), .C(n3137), .D(n32988), .Y(n32778) );
  AOI22X1 U21866 ( .A(n3233), .B(n25491), .C(n3191), .D(n23470), .Y(n32781) );
  OAI21X1 U21867 ( .A(n25404), .B(n32782), .C(n21883), .Y(n32786) );
  AOI22X1 U21868 ( .A(n3221), .B(n23307), .C(n3215), .D(n23306), .Y(n32784) );
  OAI21X1 U21869 ( .A(n25443), .B(n32912), .C(n21884), .Y(n32785) );
  NOR3X1 U21870 ( .A(n32786), .B(n22934), .C(n32785), .Y(n32797) );
  AOI22X1 U21871 ( .A(n3149), .B(n32882), .C(n3143), .D(n27218), .Y(n32789) );
  AOI22X1 U21872 ( .A(n3173), .B(n32871), .C(n3167), .D(n32877), .Y(n32787) );
  AOI22X1 U21873 ( .A(n3125), .B(n27219), .C(n3107), .D(n27217), .Y(n32790) );
  OAI21X1 U21874 ( .A(n26811), .B(n32791), .C(n21885), .Y(n32795) );
  AOI22X1 U21875 ( .A(n3131), .B(n27220), .C(n3119), .D(n27216), .Y(n32793) );
  OAI21X1 U21876 ( .A(n27115), .B(n32848), .C(n21886), .Y(n32794) );
  NOR3X1 U21877 ( .A(n22906), .B(n32795), .C(n32794), .Y(n32796) );
  NAND3X1 U21878 ( .A(n32800), .B(n32799), .C(n32798), .Y(n32801) );
  AOI22X1 U21879 ( .A(n33875), .B(n3111), .C(n33900), .D(n3105), .Y(n32802) );
  AOI22X1 U21880 ( .A(n33216), .B(n3271), .C(n33247), .D(n3265), .Y(n32804) );
  OAI21X1 U21881 ( .A(n32805), .B(n21375), .C(n21887), .Y(n32806) );
  AOI22X1 U21882 ( .A(n33806), .B(n3129), .C(n25675), .D(n3123), .Y(n32808) );
  OAI21X1 U21883 ( .A(n32809), .B(n27199), .C(n21888), .Y(n32813) );
  AOI22X1 U21884 ( .A(n26077), .B(n3147), .C(n33762), .D(n3141), .Y(n32810) );
  OAI21X1 U21885 ( .A(n32811), .B(n21378), .C(n21889), .Y(n32812) );
  NOR3X1 U21886 ( .A(n32812), .B(n32813), .C(n32814), .Y(n32845) );
  AOI22X1 U21887 ( .A(n25628), .B(n3199), .C(n33560), .D(n3193), .Y(n32817) );
  AOI22X1 U21888 ( .A(n33912), .B(n3223), .C(n33471), .D(n3217), .Y(n32815) );
  NAND3X1 U21889 ( .A(n22524), .B(n24591), .C(n24792), .Y(n32823) );
  AOI22X1 U21890 ( .A(n33399), .B(n3235), .C(n33430), .D(n3229), .Y(n32818) );
  OAI21X1 U21891 ( .A(n32980), .B(n25452), .C(n21890), .Y(n32822) );
  AOI22X1 U21892 ( .A(n33308), .B(n3253), .C(n33339), .D(n3247), .Y(n32819) );
  OAI21X1 U21893 ( .A(n32820), .B(n25453), .C(n21891), .Y(n32821) );
  AOI22X1 U21894 ( .A(n33429), .B(n3225), .C(n33462), .D(n3219), .Y(n32826) );
  AOI22X1 U21895 ( .A(n25680), .B(n3243), .C(n25657), .D(n3237), .Y(n32824) );
  AOI22X1 U21896 ( .A(n25658), .B(n3261), .C(n33295), .D(n3255), .Y(n32827) );
  OAI21X1 U21897 ( .A(n33394), .B(n21384), .C(n21892), .Y(n32830) );
  AOI22X1 U21898 ( .A(n23457), .B(RO[177]), .C(n34222), .D(n3273), .Y(n32828)
         );
  OAI21X1 U21899 ( .A(n33211), .B(n21387), .C(n21893), .Y(n32829) );
  NOR3X1 U21900 ( .A(n32829), .B(n32830), .C(n22930), .Y(n32842) );
  AOI22X1 U21901 ( .A(n33696), .B(n3159), .C(n33718), .D(n3153), .Y(n32834) );
  AOI22X1 U21902 ( .A(n21232), .B(n3177), .C(n33653), .D(n3171), .Y(n32832) );
  AOI22X1 U21903 ( .A(n33551), .B(n3195), .C(n33587), .D(n3189), .Y(n32835) );
  OAI21X1 U21904 ( .A(n32952), .B(n27207), .C(n21894), .Y(n32839) );
  AOI22X1 U21905 ( .A(n33485), .B(n3213), .C(n33508), .D(n3207), .Y(n32836) );
  OAI21X1 U21906 ( .A(n32837), .B(n25457), .C(n21895), .Y(n32838) );
  NOR3X1 U21907 ( .A(n32840), .B(n32839), .C(n32838), .Y(n32841) );
  NAND3X1 U21908 ( .A(n32845), .B(n22671), .C(n32843), .Y(n32846) );
  AOI22X1 U21909 ( .A(n3155), .B(n29836), .C(n3149), .D(n29824), .Y(n32847) );
  OAI21X1 U21910 ( .A(n27203), .B(n32848), .C(n21896), .Y(n32852) );
  AOI22X1 U21911 ( .A(n3137), .B(n29803), .C(n3131), .D(n29794), .Y(n32849) );
  OAI21X1 U21912 ( .A(n27026), .B(n32850), .C(n21897), .Y(n32851) );
  OR2X2 U21913 ( .A(n32852), .B(n32851), .Y(n32858) );
  OAI21X1 U21914 ( .A(n27120), .B(n32853), .C(n27140), .Y(n32857) );
  OAI21X1 U21915 ( .A(n27023), .B(n32854), .C(n27042), .Y(n32856) );
  NOR3X1 U21916 ( .A(n32858), .B(n32857), .C(n32856), .Y(n32891) );
  AOI22X1 U21917 ( .A(n3243), .B(n32477), .C(n3255), .D(n32478), .Y(n32861) );
  AOI22X1 U21918 ( .A(n3267), .B(n23453), .C(n3225), .D(n32480), .Y(n32859) );
  AOI22X1 U21919 ( .A(n3119), .B(n29190), .C(n3249), .D(n32957), .Y(n32862) );
  OAI21X1 U21920 ( .A(n25445), .B(n33364), .C(n21898), .Y(n32866) );
  AOI22X1 U21921 ( .A(n3107), .B(n33884), .C(RO[177]), .D(n27250), .Y(n32864)
         );
  OAI21X1 U21922 ( .A(n27189), .B(n34225), .C(n21899), .Y(n32865) );
  NOR3X1 U21923 ( .A(n22910), .B(n32866), .C(n32865), .Y(n32890) );
  AOI22X1 U21924 ( .A(n27225), .B(n3177), .C(n3189), .D(n23470), .Y(n32869) );
  AOI22X1 U21925 ( .A(n3201), .B(n32490), .C(n27298), .D(RO[179]), .Y(n32867)
         );
  AOI22X1 U21926 ( .A(n3231), .B(n25491), .C(n3183), .D(n32783), .Y(n32870) );
  OAI21X1 U21927 ( .A(n32872), .B(n27078), .C(n21900), .Y(n32876) );
  AOI22X1 U21928 ( .A(n3219), .B(n23307), .C(n3213), .D(n23306), .Y(n32873) );
  OAI21X1 U21929 ( .A(n21222), .B(n32874), .C(n21901), .Y(n32875) );
  NOR3X1 U21930 ( .A(n22914), .B(n32876), .C(n32875), .Y(n32888) );
  AOI22X1 U21931 ( .A(n32988), .B(n3135), .C(n27218), .D(n3141), .Y(n32880) );
  AOI22X1 U21932 ( .A(n27232), .B(n3159), .C(n21220), .D(n3165), .Y(n32878) );
  AOI22X1 U21933 ( .A(n27219), .B(n3123), .C(n27217), .D(n3105), .Y(n32881) );
  OAI21X1 U21934 ( .A(n32883), .B(n26996), .C(n21902), .Y(n32886) );
  OAI21X1 U21935 ( .A(n32942), .B(n27115), .C(n32884), .Y(n32885) );
  NOR3X1 U21936 ( .A(n32885), .B(n32886), .C(n22975), .Y(n32887) );
  AND2X2 U21937 ( .A(n32887), .B(n32888), .Y(n32889) );
  NAND3X1 U21938 ( .A(n32891), .B(n32890), .C(n32889), .Y(n32892) );
  AOI22X1 U21939 ( .A(n33875), .B(n3109), .C(n33900), .D(n3103), .Y(n32893) );
  OAI21X1 U21940 ( .A(n26269), .B(n32894), .C(n21903), .Y(n32899) );
  AOI22X1 U21941 ( .A(n3269), .B(n33216), .C(n3263), .D(n33247), .Y(n32896) );
  OAI21X1 U21942 ( .A(n32897), .B(n21375), .C(n21904), .Y(n32898) );
  OR2X2 U21943 ( .A(n32899), .B(n32898), .Y(n32904) );
  AOI22X1 U21944 ( .A(n33806), .B(n3127), .C(n33829), .D(n3121), .Y(n32900) );
  OAI21X1 U21945 ( .A(n27198), .B(n32901), .C(n21905), .Y(n32903) );
  OAI21X1 U21946 ( .A(n32987), .B(n21378), .C(n27143), .Y(n32902) );
  NOR3X1 U21947 ( .A(n32902), .B(n32903), .C(n32904), .Y(n32939) );
  AOI22X1 U21948 ( .A(n3197), .B(n25628), .C(n3191), .D(n33560), .Y(n32907) );
  AOI22X1 U21949 ( .A(n3221), .B(n33912), .C(n3215), .D(n33471), .Y(n32905) );
  NAND3X1 U21950 ( .A(n22527), .B(n23640), .C(n24794), .Y(n32916) );
  AOI22X1 U21951 ( .A(n3233), .B(n33399), .C(n3227), .D(n33430), .Y(n32908) );
  OAI21X1 U21952 ( .A(n25452), .B(n32909), .C(n23778), .Y(n32915) );
  AOI22X1 U21953 ( .A(n3251), .B(n33308), .C(n3245), .D(n33339), .Y(n32911) );
  OAI21X1 U21954 ( .A(n25454), .B(n32912), .C(n21906), .Y(n32914) );
  NOR3X1 U21955 ( .A(n22918), .B(n32915), .C(n32914), .Y(n32938) );
  AOI22X1 U21956 ( .A(n33429), .B(n3223), .C(n33462), .D(n3217), .Y(n32919) );
  AOI22X1 U21957 ( .A(n25680), .B(n3241), .C(n25657), .D(n3235), .Y(n32917) );
  NAND3X1 U21958 ( .A(n24126), .B(n21511), .C(n22751), .Y(n32925) );
  AOI22X1 U21959 ( .A(n25658), .B(n3259), .C(n33295), .D(n3253), .Y(n32920) );
  OAI21X1 U21960 ( .A(n32963), .B(n21384), .C(n21907), .Y(n32924) );
  AOI22X1 U21961 ( .A(n23457), .B(RO[175]), .C(n34222), .D(n3271), .Y(n32921)
         );
  OAI21X1 U21962 ( .A(n32922), .B(n21387), .C(n21908), .Y(n32923) );
  NOR3X1 U21963 ( .A(n32923), .B(n32924), .C(n22919), .Y(n32936) );
  AOI22X1 U21964 ( .A(n33696), .B(n3157), .C(n33718), .D(n3151), .Y(n32928) );
  AOI22X1 U21965 ( .A(n21232), .B(n3175), .C(n33653), .D(n3169), .Y(n32926) );
  AOI22X1 U21966 ( .A(n33551), .B(n3193), .C(n33587), .D(n3187), .Y(n32929) );
  OAI21X1 U21967 ( .A(n32977), .B(n27207), .C(n21909), .Y(n32933) );
  AOI22X1 U21968 ( .A(n33485), .B(n3211), .C(n33508), .D(n3205), .Y(n32930) );
  OAI21X1 U21969 ( .A(n32931), .B(n25455), .C(n23779), .Y(n32932) );
  NOR3X1 U21970 ( .A(n22931), .B(n32933), .C(n32932), .Y(n32935) );
  NAND3X1 U21971 ( .A(n32939), .B(n32938), .C(n32937), .Y(n32940) );
  AOI22X1 U21972 ( .A(n3147), .B(n29824), .C(n3135), .D(n25769), .Y(n32941) );
  OAI21X1 U21973 ( .A(n27205), .B(n32942), .C(n21910), .Y(n32947) );
  AOI22X1 U21974 ( .A(n3117), .B(n29190), .C(n3129), .D(n29794), .Y(n32943) );
  OAI21X1 U21975 ( .A(n27027), .B(n32944), .C(n21911), .Y(n32946) );
  AOI22X1 U21976 ( .A(n3159), .B(n23469), .C(n3153), .D(n23468), .Y(n32948) );
  OAI21X1 U21977 ( .A(n27120), .B(n32949), .C(n21912), .Y(n32955) );
  AOI22X1 U21978 ( .A(n3177), .B(n26518), .C(n3171), .D(n33639), .Y(n32951) );
  OAI21X1 U21979 ( .A(n32953), .B(n32952), .C(n23780), .Y(n32954) );
  NOR3X1 U21980 ( .A(n32954), .B(n32955), .C(n32956), .Y(n32999) );
  AOI22X1 U21981 ( .A(n3241), .B(n32477), .C(n3253), .D(n32478), .Y(n32960) );
  AOI22X1 U21982 ( .A(n3259), .B(n23451), .C(n3223), .D(n32480), .Y(n32958) );
  AOI22X1 U21983 ( .A(n3265), .B(n23452), .C(n3235), .D(n32961), .Y(n32962) );
  OAI21X1 U21984 ( .A(n32964), .B(n32963), .C(n21913), .Y(n32969) );
  AOI22X1 U21985 ( .A(n3105), .B(n33884), .C(RO[175]), .D(n27250), .Y(n32965)
         );
  OAI21X1 U21986 ( .A(n27189), .B(n32966), .C(n21914), .Y(n32968) );
  NOR3X1 U21987 ( .A(n22920), .B(n32969), .C(n32968), .Y(n32998) );
  AOI22X1 U21988 ( .A(n3175), .B(n27225), .C(n3187), .D(n23470), .Y(n32975) );
  AOI22X1 U21989 ( .A(n3193), .B(n32973), .C(n21396), .D(n29933), .Y(n32974)
         );
  AOI22X1 U21990 ( .A(n3199), .B(n32490), .C(n3169), .D(n21152), .Y(n32976) );
  OAI21X1 U21991 ( .A(n26870), .B(n32977), .C(n21915), .Y(n32982) );
  AOI22X1 U21992 ( .A(n3217), .B(n23307), .C(n3211), .D(n23306), .Y(n32979) );
  OAI21X1 U21993 ( .A(n21222), .B(n32980), .C(n21916), .Y(n32981) );
  NOR3X1 U21994 ( .A(n22924), .B(n32982), .C(n32981), .Y(n32996) );
  AOI22X1 U21995 ( .A(n3127), .B(n27220), .C(n3139), .D(n27218), .Y(n32985) );
  AOI22X1 U21996 ( .A(n3145), .B(n32882), .C(n3157), .D(n27232), .Y(n32983) );
  NAND3X1 U21997 ( .A(n22530), .B(n22732), .C(n22752), .Y(n32994) );
  AOI22X1 U21998 ( .A(n3121), .B(n27219), .C(n3103), .D(n27217), .Y(n32986) );
  OAI21X1 U21999 ( .A(n26931), .B(n32987), .C(n21917), .Y(n32993) );
  AOI22X1 U22000 ( .A(RO[177]), .B(n27298), .C(n3115), .D(n27216), .Y(n32989)
         );
  OAI21X1 U22001 ( .A(n27115), .B(n32990), .C(n21918), .Y(n32992) );
  NOR3X1 U22002 ( .A(n32993), .B(n24891), .C(n32992), .Y(n32995) );
  NAND3X1 U22003 ( .A(n32999), .B(n32997), .C(n32998), .Y(n33000) );
  AOI22X1 U22004 ( .A(n3113), .B(n33852), .C(n33875), .D(n3107), .Y(n33001) );
  OAI21X1 U22005 ( .A(n25442), .B(n33303), .C(n21919), .Y(n33006) );
  AOI22X1 U22006 ( .A(n3261), .B(n33247), .C(n3255), .D(n33277), .Y(n33003) );
  OAI21X1 U22007 ( .A(n27200), .B(n34225), .C(n21920), .Y(n33005) );
  AOI22X1 U22008 ( .A(n3125), .B(n33806), .C(n3119), .D(n33829), .Y(n33007) );
  OAI21X1 U22009 ( .A(n27195), .B(n33211), .C(n23434), .Y(n33012) );
  AOI22X1 U22010 ( .A(n3143), .B(n26077), .C(n3137), .D(n33762), .Y(n33009) );
  OAI21X1 U22011 ( .A(n21378), .B(n33010), .C(n21921), .Y(n33011) );
  NOR3X1 U22012 ( .A(n33011), .B(n33012), .C(n33013), .Y(n33048) );
  AOI22X1 U22013 ( .A(n3195), .B(n25628), .C(n3189), .D(n33560), .Y(n33016) );
  AOI22X1 U22014 ( .A(n3213), .B(n33471), .C(n3201), .D(n33517), .Y(n33014) );
  NAND3X1 U22015 ( .A(n21180), .B(n24592), .C(n24795), .Y(n33024) );
  AOI22X1 U22016 ( .A(n3225), .B(n33430), .C(n3219), .D(n33912), .Y(n33017) );
  OAI21X1 U22017 ( .A(n26078), .B(n33018), .C(n23781), .Y(n33023) );
  AOI22X1 U22018 ( .A(n3243), .B(n33339), .C(n3237), .D(n33369), .Y(n33020) );
  OAI21X1 U22019 ( .A(n21435), .B(n33394), .C(n23782), .Y(n33022) );
  NOR3X1 U22020 ( .A(n22927), .B(n33023), .C(n33022), .Y(n33047) );
  AOI22X1 U22021 ( .A(n3221), .B(n33429), .C(n3215), .D(n33462), .Y(n33027) );
  AOI22X1 U22022 ( .A(n3257), .B(n25658), .C(n3251), .D(n33295), .Y(n33028) );
  OAI21X1 U22023 ( .A(n21384), .B(n33029), .C(n21922), .Y(n33033) );
  AOI22X1 U22024 ( .A(n3275), .B(n23457), .C(n3269), .D(n34222), .Y(n33030) );
  OAI21X1 U22025 ( .A(n21387), .B(n33031), .C(n21923), .Y(n33032) );
  AOI22X1 U22026 ( .A(n3155), .B(n33696), .C(n3149), .D(n33718), .Y(n33036) );
  AOI22X1 U22027 ( .A(n3173), .B(n21232), .C(n3167), .D(n33653), .Y(n33034) );
  AOI22X1 U22028 ( .A(n3191), .B(n33551), .C(n3185), .D(n33587), .Y(n33037) );
  OAI21X1 U22029 ( .A(n27207), .B(n33038), .C(n23783), .Y(n33042) );
  AOI22X1 U22030 ( .A(n3209), .B(n33485), .C(n3203), .D(n33508), .Y(n33039) );
  OAI21X1 U22031 ( .A(n25455), .B(n33040), .C(n23784), .Y(n33041) );
  NOR3X1 U22032 ( .A(n22932), .B(n33042), .C(n33041), .Y(n33044) );
  NAND3X1 U22033 ( .A(n27902), .B(n27251), .C(n21426), .Y(n33075) );
  XOR2X1 U22034 ( .A(n22967), .B(n25611), .Y(n33059) );
  NAND3X1 U22035 ( .A(n21138), .B(n33059), .C(n34360), .Y(n33155) );
  OAI21X1 U22036 ( .A(n21154), .B(n33060), .C(T[3]), .Y(n33156) );
  XOR2X1 U22037 ( .A(n29422), .B(n33062), .Y(n33065) );
  NOR3X1 U22038 ( .A(n34441), .B(n25688), .C(n21229), .Y(n33063) );
  NAND3X1 U22039 ( .A(n27251), .B(n34443), .C(n33063), .Y(n33064) );
  AOI21X1 U22040 ( .A(n33073), .B(n33072), .C(n33086), .Y(n33070) );
  OAI21X1 U22041 ( .A(n27911), .B(n23094), .C(n27915), .Y(n33067) );
  OAI21X1 U22042 ( .A(n21154), .B(n22967), .C(n33067), .Y(n33069) );
  OAI21X1 U22043 ( .A(n34385), .B(n33069), .C(n21992), .Y(n33091) );
  OAI21X1 U22044 ( .A(n22684), .B(n33091), .C(n21992), .Y(n33071) );
  NAND3X1 U22045 ( .A(n33076), .B(n25611), .C(n21138), .Y(n33081) );
  XOR2X1 U22046 ( .A(n26072), .B(n34355), .Y(n33078) );
  FAX1 U22047 ( .A(n25619), .B(T[4]), .C(n26072), .YC(), .YS(n33080) );
  AOI21X1 U22048 ( .A(n33099), .B(n33080), .C(n33096), .Y(n33083) );
  OAI21X1 U22049 ( .A(n33082), .B(n34351), .C(n33104), .Y(n33097) );
  OAI21X1 U22050 ( .A(n33154), .B(n33158), .C(n25832), .Y(n33084) );
  OAI21X1 U22051 ( .A(n25162), .B(n25826), .C(n33084), .Y(n33144) );
  OAI21X1 U22052 ( .A(n24282), .B(n33086), .C(n23069), .Y(n33088) );
  XOR2X1 U22053 ( .A(n33088), .B(n33087), .Y(n33094) );
  NAND3X1 U22054 ( .A(n25070), .B(n33091), .C(n24872), .Y(n33093) );
  MUX2X1 U22055 ( .B(n33094), .A(n24317), .S(n33092), .Y(n33106) );
  OAI21X1 U22056 ( .A(n33096), .B(n33156), .C(n25112), .Y(n33103) );
  AOI21X1 U22057 ( .A(n33099), .B(n25112), .C(n22273), .Y(n33101) );
  MUX2X1 U22058 ( .B(n21517), .A(n22725), .S(n33100), .Y(n33105) );
  NAND3X1 U22059 ( .A(n25730), .B(n33104), .C(n33103), .Y(n33167) );
  OAI21X1 U22060 ( .A(n23099), .B(n25400), .C(n24974), .Y(n33108) );
  AOI21X1 U22061 ( .A(n25400), .B(n21230), .C(n33108), .Y(n33150) );
  AOI21X1 U22062 ( .A(n25845), .B(n25206), .C(n33110), .Y(n33109) );
  OAI21X1 U22063 ( .A(n34385), .B(n25831), .C(n21411), .Y(n33123) );
  OAI21X1 U22064 ( .A(n23139), .B(n33123), .C(n21363), .Y(n33113) );
  OAI21X1 U22065 ( .A(n23093), .B(n33110), .C(n25196), .Y(n33121) );
  NAND3X1 U22066 ( .A(n21363), .B(n25690), .C(n33121), .Y(n34255) );
  XOR2X1 U22067 ( .A(n25340), .B(n33114), .Y(n33118) );
  XOR2X1 U22068 ( .A(n25418), .B(n33114), .Y(n33117) );
  XOR2X1 U22069 ( .A(n34441), .B(T[5]), .Y(n33133) );
  OAI21X1 U22070 ( .A(n25418), .B(n23097), .C(n25337), .Y(n33116) );
  AOI22X1 U22071 ( .A(n20969), .B(n34351), .C(n33131), .D(n33116), .Y(n33137)
         );
  MUX2X1 U22072 ( .B(n33118), .A(n33117), .S(n23188), .Y(n33151) );
  OAI21X1 U22073 ( .A(n34305), .B(n25396), .C(n33151), .Y(n33119) );
  OAI21X1 U22074 ( .A(n33120), .B(n25759), .C(n33119), .Y(n33147) );
  XNOR2X1 U22075 ( .A(n33123), .B(n33121), .Y(n33127) );
  NAND3X1 U22076 ( .A(n24985), .B(n33123), .C(n22879), .Y(n33126) );
  MUX2X1 U22077 ( .B(n33127), .A(n25131), .S(n33125), .Y(n34309) );
  OAI21X1 U22078 ( .A(n33129), .B(n25340), .C(n22991), .Y(n33130) );
  AOI21X1 U22079 ( .A(n33132), .B(n22991), .C(n21522), .Y(n33138) );
  MUX2X1 U22080 ( .B(n21520), .A(n24318), .S(n23188), .Y(n33140) );
  AOI22X1 U22081 ( .A(n33142), .B(n24315), .C(n34309), .D(n33148), .Y(n33143)
         );
  AOI21X1 U22082 ( .A(n33166), .B(n26053), .C(n34434), .Y(n33149) );
  FAX1 U22083 ( .A(n33148), .B(n34323), .C(n25828), .YC(), .YS(n34420) );
  AOI22X1 U22084 ( .A(n24327), .B(n22722), .C(n27233), .D(n25862), .Y(n33173)
         );
  FAX1 U22085 ( .A(n33153), .B(n25759), .C(n25396), .YC(), .YS(n34407) );
  FAX1 U22086 ( .A(n25756), .B(n33158), .C(n33154), .YC(), .YS(n33163) );
  NAND3X1 U22087 ( .A(n25329), .B(n33156), .C(n23426), .Y(n33159) );
  XOR2X1 U22088 ( .A(n25446), .B(n33157), .Y(n34326) );
  AOI21X1 U22089 ( .A(n24259), .B(n33158), .C(n34326), .Y(n33160) );
  OAI21X1 U22090 ( .A(n34414), .B(n33161), .C(n23881), .Y(n33162) );
  OAI21X1 U22091 ( .A(n25858), .B(n33163), .C(n33162), .Y(n33164) );
  OAI21X1 U22092 ( .A(n25862), .B(n27233), .C(n33164), .Y(n33172) );
  NAND3X1 U22093 ( .A(n3773), .B(n3774), .C(n34280), .Y(n33176) );
  AOI21X1 U22094 ( .A(n33172), .B(n22678), .C(n33171), .Y(n11045) );
  NAND2X1 U22095 ( .A(n22635), .B(n23443), .Y(n33174) );
  NAND3X1 U22096 ( .A(n3774), .B(n34230), .C(n34280), .Y(n34313) );
  AOI21X1 U22097 ( .A(n22680), .B(n24249), .C(reset), .Y(n34283) );
  AOI21X1 U22098 ( .A(n22681), .B(n24250), .C(reset), .Y(n34282) );
  AOI22X1 U22099 ( .A(net95147), .B(net150130), .C(n21007), .D(net114546), .Y(
        n33181) );
  OR2X2 U22100 ( .A(reset), .B(n22122), .Y(n33885) );
  MUX2X1 U22101 ( .B(n22689), .A(n29343), .S(n34342), .Y(n33183) );
  AOI21X1 U22102 ( .A(n29400), .B(n34222), .C(n33183), .Y(n33184) );
  OAI21X1 U22103 ( .A(n33185), .B(n29211), .C(n21971), .Y(n33186) );
  AOI22X1 U22104 ( .A(n33188), .B(n33187), .C(n33188), .D(net96588), .Y(n34444) );
  AOI21X1 U22105 ( .A(n22682), .B(n24251), .C(reset), .Y(n34341) );
  AOI22X1 U22106 ( .A(n29408), .B(n33216), .C(n29425), .D(n3271), .Y(n33195)
         );
  AOI22X1 U22107 ( .A(n21219), .B(net105814), .C(n23611), .D(net114546), .Y(
        n33191) );
  OR2X2 U22108 ( .A(reset), .B(n22126), .Y(n34219) );
  AOI21X1 U22109 ( .A(n22683), .B(n24252), .C(reset), .Y(n34343) );
  AOI22X1 U22110 ( .A(n23308), .B(n29362), .C(n29414), .D(n34222), .Y(n33194)
         );
  AOI22X1 U22111 ( .A(n27292), .B(n33196), .C(n27292), .D(net96582), .Y(n34461) );
  AOI22X1 U22112 ( .A(n29386), .B(n34222), .C(n23308), .D(n29349), .Y(n33198)
         );
  AOI22X1 U22113 ( .A(n29431), .B(n3270), .C(n29398), .D(n33216), .Y(n33197)
         );
  AND2X2 U22114 ( .A(n23545), .B(n23712), .Y(n33200) );
  AOI22X1 U22115 ( .A(n33200), .B(n33199), .C(n33200), .D(net96584), .Y(n34462) );
  AOI22X1 U22116 ( .A(n23308), .B(n29408), .C(n29424), .D(n3269), .Y(n33202)
         );
  AOI22X1 U22117 ( .A(n29360), .B(n34222), .C(n29414), .D(n33216), .Y(n33201)
         );
  AOI22X1 U22118 ( .A(n27293), .B(n33203), .C(n27293), .D(net96586), .Y(n34463) );
  AOI22X1 U22119 ( .A(n29386), .B(n33216), .C(n29349), .D(n34222), .Y(n33205)
         );
  AOI22X1 U22120 ( .A(n29431), .B(n3268), .C(n23308), .D(n29400), .Y(n33204)
         );
  AND2X2 U22121 ( .A(n23549), .B(n23713), .Y(n33207) );
  AOI22X1 U22122 ( .A(n33207), .B(n33206), .C(n33207), .D(net96588), .Y(n34464) );
  MUX2X1 U22123 ( .B(n22690), .A(n29355), .S(n33216), .Y(n33209) );
  AOI21X1 U22124 ( .A(n29409), .B(n33234), .C(n33209), .Y(n33210) );
  OAI21X1 U22125 ( .A(n33211), .B(n29211), .C(n21972), .Y(n33212) );
  AOI22X1 U22126 ( .A(n33214), .B(n33213), .C(n33214), .D(net96588), .Y(n34445) );
  MUX2X1 U22127 ( .B(n22691), .A(n29343), .S(n33216), .Y(n33218) );
  AOI21X1 U22128 ( .A(n29400), .B(n33234), .C(n33218), .Y(n33219) );
  OAI21X1 U22129 ( .A(n33220), .B(n29211), .C(n21973), .Y(n33221) );
  AOI22X1 U22130 ( .A(n33223), .B(n33222), .C(n33223), .D(net96588), .Y(n34446) );
  AOI22X1 U22131 ( .A(n29409), .B(n33247), .C(n29424), .D(n3265), .Y(n33225)
         );
  AOI22X1 U22132 ( .A(n30612), .B(n29361), .C(n29414), .D(n33234), .Y(n33224)
         );
  AOI22X1 U22133 ( .A(n27284), .B(n33226), .C(n27284), .D(net96588), .Y(n34465) );
  AOI22X1 U22134 ( .A(n29386), .B(n33234), .C(n30612), .D(n29348), .Y(n33228)
         );
  AOI22X1 U22135 ( .A(n29431), .B(n3264), .C(n29397), .D(n33247), .Y(n33227)
         );
  AND2X2 U22136 ( .A(n23551), .B(n23715), .Y(n33230) );
  AOI22X1 U22137 ( .A(n33230), .B(n33229), .C(n33230), .D(net96588), .Y(n34466) );
  AOI22X1 U22138 ( .A(n30612), .B(n29409), .C(n29424), .D(n3263), .Y(n33232)
         );
  AOI22X1 U22139 ( .A(n29361), .B(n33234), .C(n29414), .D(n33247), .Y(n33231)
         );
  AOI22X1 U22140 ( .A(n27287), .B(n33233), .C(n27287), .D(net96588), .Y(n34467) );
  AOI22X1 U22141 ( .A(n29386), .B(n33247), .C(n29351), .D(n33234), .Y(n33236)
         );
  AOI22X1 U22142 ( .A(n29431), .B(n3262), .C(n30612), .D(n29399), .Y(n33235)
         );
  AND2X2 U22143 ( .A(n23554), .B(n23716), .Y(n33238) );
  AOI22X1 U22144 ( .A(n33238), .B(n33237), .C(n33238), .D(net96588), .Y(n34468) );
  MUX2X1 U22145 ( .B(n22692), .A(n29354), .S(n33247), .Y(n33240) );
  AOI21X1 U22146 ( .A(n29409), .B(n25658), .C(n33240), .Y(n33241) );
  OAI21X1 U22147 ( .A(n33242), .B(n29211), .C(n21974), .Y(n33243) );
  AOI22X1 U22148 ( .A(n33245), .B(n33244), .C(n33245), .D(net96588), .Y(n34447) );
  MUX2X1 U22149 ( .B(n22693), .A(n29343), .S(n33247), .Y(n33249) );
  AOI21X1 U22150 ( .A(n29400), .B(n25658), .C(n33249), .Y(n33250) );
  OAI21X1 U22151 ( .A(n33251), .B(n29211), .C(n21975), .Y(n33252) );
  AOI22X1 U22152 ( .A(n33254), .B(n33253), .C(n33254), .D(net96588), .Y(n34448) );
  AOI22X1 U22153 ( .A(n29409), .B(n33277), .C(n29424), .D(n3259), .Y(n33256)
         );
  AOI22X1 U22154 ( .A(n30607), .B(n29361), .C(n29414), .D(n25658), .Y(n33255)
         );
  AOI22X1 U22155 ( .A(n27277), .B(n33257), .C(n27277), .D(net96588), .Y(n34469) );
  AOI22X1 U22156 ( .A(n29386), .B(n25658), .C(n30607), .D(n29348), .Y(n33259)
         );
  AOI22X1 U22157 ( .A(n29431), .B(n21179), .C(n29398), .D(n33277), .Y(n33258)
         );
  AND2X2 U22158 ( .A(n23557), .B(n23718), .Y(n33261) );
  AOI22X1 U22159 ( .A(n33261), .B(n33260), .C(n33261), .D(net96588), .Y(n34470) );
  AOI22X1 U22160 ( .A(n30607), .B(n29409), .C(n29424), .D(n3257), .Y(n33263)
         );
  AOI22X1 U22161 ( .A(n29361), .B(n25658), .C(n29414), .D(n33277), .Y(n33262)
         );
  AOI22X1 U22162 ( .A(n27278), .B(n33264), .C(n27278), .D(net96588), .Y(n34471) );
  AOI22X1 U22163 ( .A(n29386), .B(n33277), .C(n29350), .D(n25658), .Y(n33266)
         );
  AOI22X1 U22164 ( .A(n29431), .B(n3256), .C(n30607), .D(n29400), .Y(n33265)
         );
  AND2X2 U22165 ( .A(n23559), .B(n23719), .Y(n33268) );
  AOI22X1 U22166 ( .A(n33268), .B(n33267), .C(n33268), .D(net96588), .Y(n34472) );
  MUX2X1 U22167 ( .B(n22694), .A(n29354), .S(n33277), .Y(n33270) );
  AOI21X1 U22168 ( .A(n29408), .B(n33295), .C(n33270), .Y(n33271) );
  OAI21X1 U22169 ( .A(n33272), .B(n29211), .C(n21976), .Y(n33273) );
  AOI22X1 U22170 ( .A(n33275), .B(n33274), .C(n33275), .D(net96588), .Y(n34449) );
  MUX2X1 U22171 ( .B(n22695), .A(n29343), .S(n33277), .Y(n33279) );
  AOI21X1 U22172 ( .A(n29400), .B(n33295), .C(n33279), .Y(n33280) );
  OAI21X1 U22173 ( .A(n33281), .B(n29211), .C(n21977), .Y(n33282) );
  AOI22X1 U22174 ( .A(n33284), .B(n33283), .C(n33284), .D(net96596), .Y(n34450) );
  AOI22X1 U22175 ( .A(n29409), .B(n33308), .C(n29424), .D(n3253), .Y(n33286)
         );
  AOI22X1 U22176 ( .A(n30602), .B(n29361), .C(n29414), .D(n33295), .Y(n33285)
         );
  AOI22X1 U22177 ( .A(n27279), .B(n33287), .C(n27279), .D(net96588), .Y(n34473) );
  AOI22X1 U22178 ( .A(n29386), .B(n33295), .C(n30602), .D(n29348), .Y(n33289)
         );
  AOI22X1 U22179 ( .A(n29431), .B(n3252), .C(n29397), .D(n33308), .Y(n33288)
         );
  AND2X2 U22180 ( .A(n23561), .B(n23721), .Y(n33291) );
  AOI22X1 U22181 ( .A(n33291), .B(n33290), .C(n33291), .D(net96588), .Y(n34474) );
  AOI22X1 U22182 ( .A(n30602), .B(n29409), .C(n29424), .D(n3251), .Y(n33293)
         );
  AOI22X1 U22183 ( .A(n29359), .B(n33295), .C(n29414), .D(n33308), .Y(n33292)
         );
  AOI22X1 U22184 ( .A(n27280), .B(n33294), .C(n27280), .D(net96588), .Y(n34475) );
  AOI22X1 U22185 ( .A(n29386), .B(n33308), .C(n29350), .D(n33295), .Y(n33297)
         );
  AOI22X1 U22186 ( .A(n29431), .B(n3250), .C(n30602), .D(n29398), .Y(n33296)
         );
  AND2X2 U22187 ( .A(n23564), .B(n23600), .Y(n33299) );
  AOI22X1 U22188 ( .A(n33299), .B(n33298), .C(n33299), .D(net96596), .Y(n34476) );
  MUX2X1 U22189 ( .B(n22696), .A(n29354), .S(n33308), .Y(n33301) );
  AOI21X1 U22190 ( .A(n29409), .B(n33326), .C(n33301), .Y(n33302) );
  OAI21X1 U22191 ( .A(n33303), .B(n29211), .C(n21978), .Y(n33304) );
  AOI22X1 U22192 ( .A(n33306), .B(n33305), .C(n33306), .D(net96588), .Y(n34451) );
  MUX2X1 U22193 ( .B(n22697), .A(n29343), .S(n33308), .Y(n33310) );
  AOI21X1 U22194 ( .A(n29400), .B(n33326), .C(n33310), .Y(n33311) );
  OAI21X1 U22195 ( .A(n33312), .B(n29211), .C(n21979), .Y(n33313) );
  AOI22X1 U22196 ( .A(n33315), .B(n33314), .C(n33315), .D(net96596), .Y(n34452) );
  AOI22X1 U22197 ( .A(n29409), .B(n33339), .C(n29425), .D(n3247), .Y(n33317)
         );
  AOI22X1 U22198 ( .A(n30597), .B(n29361), .C(n29414), .D(n33326), .Y(n33316)
         );
  AOI22X1 U22199 ( .A(n27285), .B(n33318), .C(n27285), .D(net96588), .Y(n34477) );
  AOI22X1 U22200 ( .A(n29386), .B(n33326), .C(n30597), .D(n29348), .Y(n33320)
         );
  AOI22X1 U22201 ( .A(n29432), .B(n3246), .C(n29397), .D(n33339), .Y(n33319)
         );
  AND2X2 U22202 ( .A(n23566), .B(n23724), .Y(n33322) );
  AOI22X1 U22203 ( .A(n33322), .B(n33321), .C(n33322), .D(net96592), .Y(n34478) );
  AOI22X1 U22204 ( .A(n30597), .B(n29409), .C(n29425), .D(n3245), .Y(n33324)
         );
  AOI22X1 U22205 ( .A(n29359), .B(n33326), .C(n29414), .D(n33339), .Y(n33323)
         );
  AOI22X1 U22206 ( .A(n27288), .B(n33325), .C(n27288), .D(net96592), .Y(n34479) );
  AOI22X1 U22207 ( .A(n29386), .B(n33339), .C(n29350), .D(n33326), .Y(n33328)
         );
  AOI22X1 U22208 ( .A(n29431), .B(n20962), .C(n30597), .D(n29396), .Y(n33327)
         );
  AND2X2 U22209 ( .A(n23568), .B(n23726), .Y(n33330) );
  AOI22X1 U22210 ( .A(n33330), .B(n33329), .C(n33330), .D(net96592), .Y(n34480) );
  MUX2X1 U22211 ( .B(n22698), .A(n29354), .S(n33339), .Y(n33332) );
  AOI21X1 U22212 ( .A(n29408), .B(n25680), .C(n33332), .Y(n33333) );
  OAI21X1 U22213 ( .A(n33334), .B(n29212), .C(n21980), .Y(n33335) );
  AOI22X1 U22214 ( .A(n33337), .B(n33336), .C(n33337), .D(net96592), .Y(n34453) );
  MUX2X1 U22215 ( .B(n22699), .A(n29344), .S(n33339), .Y(n33341) );
  AOI21X1 U22216 ( .A(n29400), .B(n25680), .C(n33341), .Y(n33342) );
  OAI21X1 U22217 ( .A(n33343), .B(n29212), .C(n21981), .Y(n33344) );
  AOI22X1 U22218 ( .A(n33346), .B(n33345), .C(n33346), .D(net96592), .Y(n34454) );
  AOI22X1 U22219 ( .A(n29408), .B(n33369), .C(n29428), .D(n3241), .Y(n33348)
         );
  AOI22X1 U22220 ( .A(n30592), .B(n29361), .C(n29414), .D(n25680), .Y(n33347)
         );
  AOI22X1 U22221 ( .A(n27286), .B(n33349), .C(n27286), .D(net96592), .Y(n34481) );
  AOI22X1 U22222 ( .A(n29386), .B(n25680), .C(n30592), .D(n29348), .Y(n33351)
         );
  AOI22X1 U22223 ( .A(n29431), .B(n3240), .C(n29397), .D(n33369), .Y(n33350)
         );
  AND2X2 U22224 ( .A(n23571), .B(n23728), .Y(n33353) );
  AOI22X1 U22225 ( .A(n33353), .B(n33352), .C(n33353), .D(net96592), .Y(n34482) );
  AOI22X1 U22226 ( .A(n30592), .B(n29409), .C(n29425), .D(n3239), .Y(n33355)
         );
  AOI22X1 U22227 ( .A(n29360), .B(n25680), .C(n29414), .D(n33369), .Y(n33354)
         );
  AOI22X1 U22228 ( .A(n27289), .B(n33356), .C(n27289), .D(net96592), .Y(n34483) );
  AOI22X1 U22229 ( .A(n29387), .B(n33369), .C(n29349), .D(n25680), .Y(n33358)
         );
  AOI22X1 U22230 ( .A(n29431), .B(n3238), .C(n30592), .D(n29399), .Y(n33357)
         );
  AND2X2 U22231 ( .A(n23574), .B(n23730), .Y(n33360) );
  AOI22X1 U22232 ( .A(n33360), .B(n33359), .C(n33360), .D(net96592), .Y(n34484) );
  MUX2X1 U22233 ( .B(n22700), .A(n29355), .S(n33369), .Y(n33362) );
  AOI21X1 U22234 ( .A(n29409), .B(n25657), .C(n33362), .Y(n33363) );
  OAI21X1 U22235 ( .A(n33364), .B(n29212), .C(n21982), .Y(n33365) );
  AOI22X1 U22236 ( .A(n33367), .B(n33366), .C(n33367), .D(net96592), .Y(n34455) );
  MUX2X1 U22237 ( .B(n22701), .A(n29344), .S(n33369), .Y(n33371) );
  AOI21X1 U22238 ( .A(n29400), .B(n25657), .C(n33371), .Y(n33372) );
  OAI21X1 U22239 ( .A(n33373), .B(n29212), .C(n23882), .Y(n33374) );
  AOI22X1 U22240 ( .A(n33376), .B(n33375), .C(n33376), .D(net96592), .Y(n34456) );
  AOI22X1 U22241 ( .A(n29408), .B(n33399), .C(n29425), .D(n3235), .Y(n33378)
         );
  AOI22X1 U22242 ( .A(n30587), .B(n29362), .C(n29414), .D(n25657), .Y(n33377)
         );
  AOI22X1 U22243 ( .A(n27290), .B(n33379), .C(n27290), .D(net96588), .Y(n34485) );
  AOI22X1 U22244 ( .A(n29386), .B(n25657), .C(n30587), .D(n29348), .Y(n33381)
         );
  AOI22X1 U22245 ( .A(n29431), .B(n3234), .C(n29397), .D(n33399), .Y(n33380)
         );
  AND2X2 U22246 ( .A(n23577), .B(n23732), .Y(n33383) );
  AOI22X1 U22247 ( .A(n33383), .B(n33382), .C(n33383), .D(net96592), .Y(n34486) );
  AOI22X1 U22248 ( .A(n30587), .B(n29409), .C(n29425), .D(n3233), .Y(n33385)
         );
  AOI22X1 U22249 ( .A(n29360), .B(n25657), .C(n29414), .D(n33399), .Y(n33384)
         );
  AOI22X1 U22250 ( .A(n29387), .B(n33399), .C(n29349), .D(n25657), .Y(n33388)
         );
  AOI22X1 U22251 ( .A(n29432), .B(n3232), .C(n30587), .D(n29396), .Y(n33387)
         );
  AND2X2 U22252 ( .A(n23581), .B(n23733), .Y(n33390) );
  AOI22X1 U22253 ( .A(n33390), .B(n33389), .C(n33390), .D(net96588), .Y(n34488) );
  MUX2X1 U22254 ( .B(n22702), .A(n29355), .S(n33399), .Y(n33392) );
  AOI21X1 U22255 ( .A(n29408), .B(n33417), .C(n33392), .Y(n33393) );
  OAI21X1 U22256 ( .A(n33394), .B(n29212), .C(n21983), .Y(n33395) );
  AOI22X1 U22257 ( .A(n33397), .B(n33396), .C(n33397), .D(net96588), .Y(n34457) );
  MUX2X1 U22258 ( .B(n22703), .A(n29344), .S(n33399), .Y(n33401) );
  AOI21X1 U22259 ( .A(n29400), .B(n33417), .C(n33401), .Y(n33402) );
  OAI21X1 U22260 ( .A(n33403), .B(n29212), .C(n21984), .Y(n33404) );
  AOI22X1 U22261 ( .A(n33406), .B(n33405), .C(n33406), .D(net96592), .Y(n34458) );
  AOI22X1 U22262 ( .A(n29408), .B(n33430), .C(n29425), .D(n3229), .Y(n33408)
         );
  AOI22X1 U22263 ( .A(n30582), .B(n29361), .C(n29414), .D(n33417), .Y(n33407)
         );
  AOI22X1 U22264 ( .A(n27282), .B(n33409), .C(n27282), .D(net96596), .Y(n34489) );
  AOI22X1 U22265 ( .A(n29387), .B(n33417), .C(n30582), .D(n29348), .Y(n33411)
         );
  AOI22X1 U22266 ( .A(n29432), .B(n3228), .C(n29397), .D(n33430), .Y(n33410)
         );
  AND2X2 U22267 ( .A(n23583), .B(n23735), .Y(n33413) );
  AOI22X1 U22268 ( .A(n33413), .B(n33412), .C(n33413), .D(net96588), .Y(n34490) );
  AOI22X1 U22269 ( .A(n30582), .B(n29409), .C(n29425), .D(n3227), .Y(n33415)
         );
  AOI22X1 U22270 ( .A(n29360), .B(n33417), .C(n29414), .D(n33430), .Y(n33414)
         );
  AOI22X1 U22271 ( .A(n27291), .B(n33416), .C(n27291), .D(net96588), .Y(n34491) );
  AOI22X1 U22272 ( .A(n29386), .B(n33430), .C(n29349), .D(n33417), .Y(n33419)
         );
  AOI22X1 U22273 ( .A(n29432), .B(n3226), .C(n30582), .D(n29396), .Y(n33418)
         );
  AND2X2 U22274 ( .A(n23585), .B(n23737), .Y(n33421) );
  AOI22X1 U22275 ( .A(n33421), .B(n33420), .C(n33421), .D(net96596), .Y(n34492) );
  MUX2X1 U22276 ( .B(n22704), .A(n29355), .S(n33430), .Y(n33423) );
  AOI21X1 U22277 ( .A(n29408), .B(n33429), .C(n33423), .Y(n33424) );
  OAI21X1 U22278 ( .A(n33425), .B(n29212), .C(n21985), .Y(n33426) );
  AOI22X1 U22279 ( .A(n33428), .B(n33427), .C(n33428), .D(net96596), .Y(n34459) );
  AOI22X1 U22280 ( .A(n29399), .B(n25774), .C(n12026), .D(net96558), .Y(n33434) );
  MUX2X1 U22281 ( .B(n22705), .A(n29344), .S(n33430), .Y(n33432) );
  AOI21X1 U22282 ( .A(n29432), .B(n3224), .C(n33432), .Y(n33433) );
  AOI22X1 U22283 ( .A(n12025), .B(net96558), .C(n29407), .D(n20856), .Y(n33437) );
  AOI22X1 U22284 ( .A(n30577), .B(n29361), .C(n29414), .D(n25774), .Y(n33435)
         );
  NAND3X1 U22285 ( .A(n22533), .B(n24593), .C(n24796), .Y(n21519) );
  AOI22X1 U22286 ( .A(n12023), .B(net96560), .C(n30577), .D(n29406), .Y(n33440) );
  AOI22X1 U22287 ( .A(n29359), .B(n33429), .C(n29414), .D(n20856), .Y(n33438)
         );
  NAND3X1 U22288 ( .A(n24797), .B(n24594), .C(n22536), .Y(n21516) );
  AOI22X1 U22289 ( .A(n12022), .B(net96558), .C(n29350), .D(n25774), .Y(n33443) );
  AOI22X1 U22290 ( .A(n30577), .B(n29400), .C(n29425), .D(n3220), .Y(n33441)
         );
  NAND3X1 U22291 ( .A(n22539), .B(n24595), .C(n24798), .Y(n21515) );
  MUX2X1 U22292 ( .B(n24284), .A(n29355), .S(n20856), .Y(n33445) );
  AOI21X1 U22293 ( .A(n12021), .B(net96574), .C(n33445), .Y(n33447) );
  AOI22X1 U22294 ( .A(n29408), .B(n33462), .C(n29425), .D(n3219), .Y(n33446)
         );
  MUX2X1 U22295 ( .B(n24285), .A(n29344), .S(n20856), .Y(n33450) );
  AOI22X1 U22296 ( .A(n29398), .B(n33462), .C(n29425), .D(n3218), .Y(n33451)
         );
  AOI22X1 U22297 ( .A(n12019), .B(net96560), .C(n29407), .D(n33471), .Y(n33455) );
  AOI22X1 U22298 ( .A(n30572), .B(n29362), .C(n29414), .D(n33462), .Y(n33453)
         );
  NAND3X1 U22299 ( .A(n24799), .B(n24596), .C(n22542), .Y(n21510) );
  AOI22X1 U22300 ( .A(n12018), .B(net96560), .C(n30572), .D(n29348), .Y(n33458) );
  AOI22X1 U22301 ( .A(n29399), .B(n33471), .C(n29425), .D(n3216), .Y(n33456)
         );
  NAND3X1 U22302 ( .A(n22545), .B(n24597), .C(n24800), .Y(n21509) );
  AOI22X1 U22303 ( .A(n12017), .B(net96560), .C(n30572), .D(n29406), .Y(n33461) );
  AOI22X1 U22304 ( .A(n29359), .B(n33462), .C(n29414), .D(n33471), .Y(n33459)
         );
  NAND3X1 U22305 ( .A(n22548), .B(n24598), .C(n24801), .Y(n21507) );
  AOI22X1 U22306 ( .A(n12016), .B(net96560), .C(n29350), .D(n33462), .Y(n33465) );
  AOI22X1 U22307 ( .A(n30572), .B(n29399), .C(n29425), .D(n3214), .Y(n33463)
         );
  NAND3X1 U22308 ( .A(n22551), .B(n24599), .C(n24802), .Y(n21506) );
  MUX2X1 U22309 ( .B(n22706), .A(n29355), .S(n33471), .Y(n33467) );
  AOI22X1 U22310 ( .A(n29408), .B(n33485), .C(n29426), .D(n3213), .Y(n33468)
         );
  MUX2X1 U22311 ( .B(n24286), .A(n29344), .S(n33471), .Y(n33473) );
  AOI22X1 U22312 ( .A(n29399), .B(n33485), .C(n29426), .D(n3212), .Y(n33474)
         );
  AOI22X1 U22313 ( .A(n12013), .B(net96560), .C(n29407), .D(n33494), .Y(n33478) );
  AOI22X1 U22314 ( .A(n30567), .B(n29362), .C(n29414), .D(n33485), .Y(n33476)
         );
  NAND3X1 U22315 ( .A(n24128), .B(n24600), .C(n22753), .Y(n21501) );
  AOI22X1 U22316 ( .A(n12012), .B(net96562), .C(n30567), .D(n29349), .Y(n33481) );
  AOI22X1 U22317 ( .A(n29399), .B(n33494), .C(n29426), .D(n3210), .Y(n33479)
         );
  NAND3X1 U22318 ( .A(n24129), .B(n24601), .C(n22754), .Y(n21500) );
  AOI22X1 U22319 ( .A(n12011), .B(net96558), .C(n30567), .D(n29405), .Y(n33484) );
  AOI22X1 U22320 ( .A(n29359), .B(n33485), .C(n29414), .D(n33494), .Y(n33482)
         );
  NAND3X1 U22321 ( .A(n24130), .B(n24602), .C(n22755), .Y(n21498) );
  AOI22X1 U22322 ( .A(n12010), .B(net96570), .C(n29350), .D(n33485), .Y(n33488) );
  AOI22X1 U22323 ( .A(n30567), .B(n29400), .C(n29426), .D(n3208), .Y(n33486)
         );
  NAND3X1 U22324 ( .A(n24131), .B(n24603), .C(n22756), .Y(n21497) );
  MUX2X1 U22325 ( .B(n24287), .A(n29355), .S(n33494), .Y(n33490) );
  AOI21X1 U22326 ( .A(n12009), .B(net96574), .C(n33490), .Y(n33492) );
  AOI22X1 U22327 ( .A(n29407), .B(n33508), .C(n29426), .D(n3207), .Y(n33491)
         );
  MUX2X1 U22328 ( .B(n24288), .A(n29344), .S(n33494), .Y(n33496) );
  AOI21X1 U22329 ( .A(n12008), .B(net96574), .C(n33496), .Y(n33498) );
  AOI22X1 U22330 ( .A(n29398), .B(n33508), .C(n29426), .D(n3206), .Y(n33497)
         );
  AOI22X1 U22331 ( .A(net96560), .B(n12007), .C(n29407), .D(n33517), .Y(n33501) );
  AOI22X1 U22332 ( .A(n23273), .B(n29362), .C(n29414), .D(n33508), .Y(n33499)
         );
  NAND3X1 U22333 ( .A(n22554), .B(n24604), .C(n24803), .Y(n21492) );
  AOI22X1 U22334 ( .A(n12006), .B(net96570), .C(n23273), .D(n29349), .Y(n33504) );
  AOI22X1 U22335 ( .A(n29398), .B(n33517), .C(n29426), .D(n3204), .Y(n33502)
         );
  NAND3X1 U22336 ( .A(n22557), .B(n24605), .C(n24804), .Y(n21491) );
  AOI22X1 U22337 ( .A(n12005), .B(net96560), .C(n23273), .D(n29406), .Y(n33507) );
  AOI22X1 U22338 ( .A(n29359), .B(n33508), .C(n29414), .D(n33517), .Y(n33505)
         );
  NAND3X1 U22339 ( .A(n22560), .B(n24606), .C(n24805), .Y(n21489) );
  AOI22X1 U22340 ( .A(n12004), .B(net96570), .C(n29351), .D(n33508), .Y(n33511) );
  AOI22X1 U22341 ( .A(n23273), .B(n29400), .C(n29426), .D(n3202), .Y(n33509)
         );
  NAND3X1 U22342 ( .A(n24132), .B(n24607), .C(n22757), .Y(n21488) );
  MUX2X1 U22343 ( .B(n22707), .A(n29355), .S(n33517), .Y(n33513) );
  AOI21X1 U22344 ( .A(n12003), .B(net96574), .C(n33513), .Y(n33515) );
  AOI22X1 U22345 ( .A(n29407), .B(n33531), .C(n29426), .D(n3201), .Y(n33514)
         );
  MUX2X1 U22346 ( .B(n24289), .A(n29344), .S(n33517), .Y(n33519) );
  AOI22X1 U22347 ( .A(n29398), .B(n33531), .C(n29426), .D(n25775), .Y(n33520)
         );
  AOI22X1 U22348 ( .A(n12001), .B(net96560), .C(n29407), .D(n33538), .Y(n33524) );
  AOI22X1 U22349 ( .A(n30558), .B(n29362), .C(n29414), .D(n33531), .Y(n33522)
         );
  NAND3X1 U22350 ( .A(n24133), .B(n24608), .C(n22758), .Y(n21483) );
  AOI22X1 U22351 ( .A(n12000), .B(net96570), .C(n30558), .D(n29349), .Y(n33527) );
  AOI22X1 U22352 ( .A(n29398), .B(n33538), .C(n29426), .D(n3198), .Y(n33525)
         );
  NAND3X1 U22353 ( .A(n24134), .B(n24609), .C(n22759), .Y(n21482) );
  AOI22X1 U22354 ( .A(n11999), .B(net96558), .C(n30558), .D(n29406), .Y(n33530) );
  AOI22X1 U22355 ( .A(n29359), .B(n33531), .C(n29414), .D(n33538), .Y(n33528)
         );
  NAND3X1 U22356 ( .A(n24135), .B(n24610), .C(n22760), .Y(n21480) );
  AOI22X1 U22357 ( .A(n11998), .B(net96570), .C(n29349), .D(n33531), .Y(n33534) );
  AOI22X1 U22358 ( .A(n30558), .B(n29400), .C(n29426), .D(n3196), .Y(n33532)
         );
  NAND3X1 U22359 ( .A(n22563), .B(n24611), .C(n24806), .Y(n21479) );
  AOI22X1 U22360 ( .A(n11997), .B(net96560), .C(n29407), .D(n33551), .Y(n33537) );
  AOI22X1 U22361 ( .A(n29360), .B(n25628), .C(n23305), .D(n29414), .Y(n33535)
         );
  NAND3X1 U22362 ( .A(n24136), .B(n24612), .C(n22761), .Y(n21477) );
  AOI22X1 U22363 ( .A(n11996), .B(net96568), .C(n29350), .D(n33538), .Y(n33541) );
  AOI22X1 U22364 ( .A(n29398), .B(n33551), .C(n29426), .D(n3194), .Y(n33539)
         );
  NAND3X1 U22365 ( .A(n24807), .B(n24613), .C(n22566), .Y(n21476) );
  AOI22X1 U22366 ( .A(n11995), .B(net96560), .C(n29407), .D(n33573), .Y(n33544) );
  AOI22X1 U22367 ( .A(n29886), .B(n29362), .C(n29414), .D(n33551), .Y(n33542)
         );
  NAND3X1 U22368 ( .A(n24137), .B(n24614), .C(n22762), .Y(n21474) );
  AOI22X1 U22369 ( .A(n11994), .B(net96564), .C(n29886), .D(n29349), .Y(n33547) );
  AOI22X1 U22370 ( .A(n29398), .B(n33573), .C(n29427), .D(n3192), .Y(n33545)
         );
  NAND3X1 U22371 ( .A(n22569), .B(n24615), .C(n24808), .Y(n21473) );
  AOI22X1 U22372 ( .A(n11993), .B(net96560), .C(n29886), .D(n29406), .Y(n33550) );
  AOI22X1 U22373 ( .A(n29360), .B(n33551), .C(n29414), .D(n33573), .Y(n33548)
         );
  NAND3X1 U22374 ( .A(n22572), .B(n24616), .C(n24809), .Y(n21471) );
  AOI22X1 U22375 ( .A(n11992), .B(net96564), .C(n29350), .D(n33551), .Y(n33554) );
  AOI22X1 U22376 ( .A(n29886), .B(n29400), .C(n29427), .D(n3190), .Y(n33552)
         );
  NAND3X1 U22377 ( .A(n22575), .B(n24617), .C(n24810), .Y(n21470) );
  AOI22X1 U22378 ( .A(n29336), .B(n33587), .C(n29332), .D(n33555), .Y(n33567)
         );
  NAND2X1 U22379 ( .A(n29341), .B(n24975), .Y(n33566) );
  NOR3X1 U22380 ( .A(n30062), .B(n14373), .C(n25597), .Y(n33564) );
  NOR3X1 U22381 ( .A(n33564), .B(n33563), .C(n33562), .Y(n33565) );
  NAND3X1 U22382 ( .A(n33567), .B(n33566), .C(n33565), .Y(n22376) );
  MUX2X1 U22383 ( .B(n22708), .A(n29355), .S(n33573), .Y(n33569) );
  AOI21X1 U22384 ( .A(n11991), .B(net96574), .C(n33569), .Y(n33571) );
  AOI22X1 U22385 ( .A(n29407), .B(n33587), .C(n29427), .D(n3189), .Y(n33570)
         );
  MUX2X1 U22386 ( .B(n24290), .A(n29344), .S(n33573), .Y(n33575) );
  AOI21X1 U22387 ( .A(n11990), .B(net96574), .C(n33575), .Y(n33577) );
  AOI22X1 U22388 ( .A(n29398), .B(n33587), .C(n29427), .D(n3188), .Y(n33576)
         );
  AOI22X1 U22389 ( .A(n11989), .B(net96560), .C(n29407), .D(n26521), .Y(n33580) );
  AOI22X1 U22390 ( .A(n23304), .B(n29362), .C(n29414), .D(n33587), .Y(n33578)
         );
  NAND3X1 U22391 ( .A(n22578), .B(n24618), .C(n24811), .Y(n21464) );
  AOI22X1 U22392 ( .A(n11988), .B(net96564), .C(n23304), .D(n29348), .Y(n33583) );
  AOI22X1 U22393 ( .A(n29398), .B(n26521), .C(n29427), .D(n3186), .Y(n33581)
         );
  NAND3X1 U22394 ( .A(n22581), .B(n24619), .C(n24812), .Y(n21463) );
  AOI22X1 U22395 ( .A(net96572), .B(n11987), .C(n23304), .D(n29406), .Y(n33586) );
  AOI22X1 U22396 ( .A(n29359), .B(n33587), .C(n29414), .D(n26521), .Y(n33584)
         );
  NAND3X1 U22397 ( .A(n22584), .B(n24620), .C(n24813), .Y(n21461) );
  AOI22X1 U22398 ( .A(n11986), .B(net96572), .C(n29350), .D(n33587), .Y(n33590) );
  AOI22X1 U22399 ( .A(n23304), .B(n29399), .C(n29427), .D(n3184), .Y(n33588)
         );
  NAND3X1 U22400 ( .A(n22587), .B(n24621), .C(n24814), .Y(n21460) );
  MUX2X1 U22401 ( .B(n22709), .A(n29355), .S(n26521), .Y(n33592) );
  AOI21X1 U22402 ( .A(n11985), .B(net96574), .C(n33592), .Y(n33594) );
  AOI22X1 U22403 ( .A(n29407), .B(n33609), .C(n29427), .D(n3183), .Y(n33593)
         );
  MUX2X1 U22404 ( .B(n24291), .A(n29344), .S(n26521), .Y(n33597) );
  AOI21X1 U22405 ( .A(n11984), .B(net96574), .C(n33597), .Y(n33599) );
  AOI22X1 U22406 ( .A(n29399), .B(n33609), .C(n29427), .D(n3182), .Y(n33598)
         );
  AOI22X1 U22407 ( .A(n11983), .B(net96572), .C(n29407), .D(n26518), .Y(n33602) );
  AOI22X1 U22408 ( .A(n30546), .B(n29362), .C(n29414), .D(n33609), .Y(n33600)
         );
  NAND3X1 U22409 ( .A(n22590), .B(n24622), .C(n24815), .Y(n21455) );
  AOI22X1 U22410 ( .A(n11982), .B(net96564), .C(n30546), .D(n29349), .Y(n33605) );
  AOI22X1 U22411 ( .A(n29398), .B(n26518), .C(n29427), .D(n3180), .Y(n33603)
         );
  NAND3X1 U22412 ( .A(n22593), .B(n24623), .C(n24816), .Y(n21454) );
  AOI22X1 U22413 ( .A(n11981), .B(net96572), .C(n30546), .D(n29406), .Y(n33608) );
  AOI22X1 U22414 ( .A(n29359), .B(n33609), .C(n29414), .D(n26518), .Y(n33606)
         );
  NAND3X1 U22415 ( .A(n22596), .B(n24624), .C(n24817), .Y(n21452) );
  AOI22X1 U22416 ( .A(n11980), .B(net96564), .C(n29351), .D(n33609), .Y(n33612) );
  AOI22X1 U22417 ( .A(n30546), .B(n29400), .C(n29427), .D(n3178), .Y(n33610)
         );
  NAND3X1 U22418 ( .A(n22599), .B(n24625), .C(n24818), .Y(n21451) );
  MUX2X1 U22419 ( .B(n22710), .A(n29355), .S(n26518), .Y(n33614) );
  AOI22X1 U22420 ( .A(n29407), .B(n21232), .C(n29427), .D(n3177), .Y(n33615)
         );
  MUX2X1 U22421 ( .B(n24292), .A(n29344), .S(n26518), .Y(n33619) );
  AOI21X1 U22422 ( .A(n11978), .B(net96572), .C(n33619), .Y(n33621) );
  AOI22X1 U22423 ( .A(n29399), .B(n21232), .C(n29427), .D(n3176), .Y(n33620)
         );
  AOI22X1 U22424 ( .A(n11977), .B(net96570), .C(n29407), .D(n33639), .Y(n33624) );
  AOI22X1 U22425 ( .A(n30541), .B(n29362), .C(n29414), .D(n21232), .Y(n33622)
         );
  NAND3X1 U22426 ( .A(n22602), .B(n24626), .C(n24819), .Y(n21446) );
  AOI22X1 U22427 ( .A(n11976), .B(net96572), .C(n30541), .D(n29349), .Y(n33627) );
  AOI22X1 U22428 ( .A(n29398), .B(n33639), .C(n29427), .D(n3174), .Y(n33625)
         );
  NAND3X1 U22429 ( .A(n22605), .B(n24627), .C(n24820), .Y(n21445) );
  AOI22X1 U22430 ( .A(n11975), .B(net96570), .C(n30541), .D(n29406), .Y(n33630) );
  AOI22X1 U22431 ( .A(n29360), .B(n21232), .C(n29414), .D(n33639), .Y(n33628)
         );
  NAND3X1 U22432 ( .A(n22608), .B(n24628), .C(n24821), .Y(n21443) );
  AOI22X1 U22433 ( .A(n11974), .B(net96572), .C(n29350), .D(n21232), .Y(n33633) );
  AOI22X1 U22434 ( .A(n30541), .B(n29400), .C(n29428), .D(n3172), .Y(n33631)
         );
  NAND3X1 U22435 ( .A(n22611), .B(n24629), .C(n24822), .Y(n21442) );
  MUX2X1 U22436 ( .B(n22711), .A(n29355), .S(n33639), .Y(n33635) );
  AOI21X1 U22437 ( .A(n11973), .B(net96572), .C(n33635), .Y(n33637) );
  AOI22X1 U22438 ( .A(n29408), .B(n33653), .C(n29428), .D(n3171), .Y(n33636)
         );
  MUX2X1 U22439 ( .B(n24293), .A(n29345), .S(n33639), .Y(n33641) );
  AOI21X1 U22440 ( .A(n11972), .B(net96572), .C(n33641), .Y(n33643) );
  AOI22X1 U22441 ( .A(n29399), .B(n33653), .C(n29428), .D(n3170), .Y(n33642)
         );
  AOI22X1 U22442 ( .A(n11971), .B(net96570), .C(n29407), .D(n26519), .Y(n33646) );
  AOI22X1 U22443 ( .A(n30536), .B(n29362), .C(n29414), .D(n33653), .Y(n33644)
         );
  NAND3X1 U22444 ( .A(n22614), .B(n24630), .C(n24823), .Y(n21437) );
  AOI22X1 U22445 ( .A(n11970), .B(net96570), .C(n30536), .D(n29348), .Y(n33649) );
  AOI22X1 U22446 ( .A(n29399), .B(n26519), .C(n29428), .D(n3168), .Y(n33647)
         );
  NAND3X1 U22447 ( .A(n22617), .B(n24631), .C(n24824), .Y(n21436) );
  AOI22X1 U22448 ( .A(n11969), .B(net96570), .C(n30536), .D(n29405), .Y(n33652) );
  AOI22X1 U22449 ( .A(n29360), .B(n33653), .C(n29414), .D(n26519), .Y(n33650)
         );
  NAND3X1 U22450 ( .A(n22620), .B(n24632), .C(n24825), .Y(n21434) );
  AOI22X1 U22451 ( .A(n11968), .B(net96562), .C(n29349), .D(n33653), .Y(n33656) );
  AOI22X1 U22452 ( .A(n30536), .B(n29399), .C(n29428), .D(n3166), .Y(n33654)
         );
  NAND3X1 U22453 ( .A(n22623), .B(n24633), .C(n24826), .Y(n21433) );
  MUX2X1 U22454 ( .B(n27047), .A(n29356), .S(n26519), .Y(n33658) );
  AOI21X1 U22455 ( .A(n11967), .B(net96572), .C(n33658), .Y(n33660) );
  AOI22X1 U22456 ( .A(n29408), .B(n33661), .C(n29428), .D(n3165), .Y(n33659)
         );
  MUX2X1 U22457 ( .B(n26964), .A(n29345), .S(n26519), .Y(n33663) );
  AOI21X1 U22458 ( .A(n11966), .B(net96572), .C(n33663), .Y(n33665) );
  AOI22X1 U22459 ( .A(n29399), .B(n33661), .C(n29428), .D(n21181), .Y(n33664)
         );
  AOI22X1 U22460 ( .A(n11965), .B(net96564), .C(n29407), .D(n23469), .Y(n33668) );
  AOI22X1 U22461 ( .A(n23303), .B(n29362), .C(n29414), .D(n33661), .Y(n33666)
         );
  NAND3X1 U22462 ( .A(n22638), .B(n24634), .C(n24827), .Y(n21428) );
  AOI22X1 U22463 ( .A(n11964), .B(net96562), .C(n23303), .D(n29348), .Y(n33671) );
  AOI22X1 U22464 ( .A(n29399), .B(n23469), .C(n29428), .D(n3162), .Y(n33669)
         );
  NAND3X1 U22465 ( .A(n22639), .B(n24635), .C(n24828), .Y(n21427) );
  AOI22X1 U22466 ( .A(n11963), .B(net96564), .C(n23303), .D(n29406), .Y(n33674) );
  AOI22X1 U22467 ( .A(n29359), .B(n33661), .C(n29414), .D(n23469), .Y(n33672)
         );
  NAND3X1 U22468 ( .A(n22640), .B(n24636), .C(n24829), .Y(n21425) );
  AOI22X1 U22469 ( .A(n29350), .B(n33661), .C(n23303), .D(n29396), .Y(n33677)
         );
  AOI22X1 U22470 ( .A(n11962), .B(net96562), .C(n29428), .D(n3160), .Y(n33675)
         );
  NAND3X1 U22471 ( .A(n24138), .B(n24637), .C(n22763), .Y(n21424) );
  AOI22X1 U22472 ( .A(n29408), .B(n33696), .C(n11961), .D(net96558), .Y(n33681) );
  MUX2X1 U22473 ( .B(n22712), .A(n29356), .S(n23469), .Y(n33679) );
  AOI21X1 U22474 ( .A(n29433), .B(n25693), .C(n33679), .Y(n33680) );
  AOI22X1 U22475 ( .A(n29399), .B(n33696), .C(n11960), .D(net96558), .Y(n33686) );
  MUX2X1 U22476 ( .B(n24294), .A(n29345), .S(n23469), .Y(n33684) );
  AOI21X1 U22477 ( .A(n29433), .B(n3158), .C(n33684), .Y(n33685) );
  AOI22X1 U22478 ( .A(n11959), .B(net96572), .C(n29407), .D(n23468), .Y(n33689) );
  AOI22X1 U22479 ( .A(n23302), .B(n29362), .C(n29414), .D(n33696), .Y(n33687)
         );
  NAND3X1 U22480 ( .A(n22641), .B(n24638), .C(n24830), .Y(n21419) );
  AOI22X1 U22481 ( .A(n23302), .B(n29351), .C(n29397), .D(n23468), .Y(n33692)
         );
  AOI22X1 U22482 ( .A(n11958), .B(net96562), .C(n29428), .D(n3156), .Y(n33690)
         );
  NAND3X1 U22483 ( .A(n24139), .B(n24639), .C(n22764), .Y(n21418) );
  AOI22X1 U22484 ( .A(n11957), .B(net96572), .C(n23302), .D(n29405), .Y(n33695) );
  AOI22X1 U22485 ( .A(n29359), .B(n33696), .C(n29414), .D(n23468), .Y(n33693)
         );
  NAND3X1 U22486 ( .A(n22642), .B(n24640), .C(n24831), .Y(n21416) );
  AOI22X1 U22487 ( .A(n29350), .B(n33696), .C(n23302), .D(n29396), .Y(n33699)
         );
  AOI22X1 U22488 ( .A(n11956), .B(net96562), .C(n29428), .D(n25776), .Y(n33697) );
  NAND3X1 U22489 ( .A(n24140), .B(n24641), .C(n22765), .Y(n21415) );
  AOI22X1 U22490 ( .A(n29408), .B(n33718), .C(n11955), .D(net96558), .Y(n33703) );
  MUX2X1 U22491 ( .B(n22713), .A(n29356), .S(n23468), .Y(n33701) );
  AOI21X1 U22492 ( .A(n29433), .B(n3153), .C(n33701), .Y(n33702) );
  MUX2X1 U22493 ( .B(n24295), .A(n29345), .S(n23468), .Y(n33706) );
  AOI21X1 U22494 ( .A(n29433), .B(n21070), .C(n33706), .Y(n33707) );
  AOI22X1 U22495 ( .A(n11953), .B(net96562), .C(n29407), .D(n26060), .Y(n33711) );
  AOI22X1 U22496 ( .A(n23300), .B(n29362), .C(n29414), .D(n33718), .Y(n33709)
         );
  NAND3X1 U22497 ( .A(n22643), .B(n24642), .C(n24832), .Y(n21410) );
  AOI22X1 U22498 ( .A(n23300), .B(n29351), .C(n29397), .D(n23467), .Y(n33714)
         );
  AOI22X1 U22499 ( .A(n11952), .B(net96562), .C(n29429), .D(n3150), .Y(n33712)
         );
  NAND3X1 U22500 ( .A(n24141), .B(n24643), .C(n22766), .Y(n21409) );
  AOI22X1 U22501 ( .A(n11951), .B(net96562), .C(n23300), .D(n29406), .Y(n33717) );
  AOI22X1 U22502 ( .A(n29359), .B(n33718), .C(n29414), .D(n26060), .Y(n33715)
         );
  NAND3X1 U22503 ( .A(n22644), .B(n24644), .C(n24833), .Y(n21407) );
  AOI22X1 U22504 ( .A(n29350), .B(n33718), .C(n23300), .D(n29396), .Y(n33721)
         );
  AOI22X1 U22505 ( .A(n11950), .B(net96562), .C(n29429), .D(n3148), .Y(n33719)
         );
  NAND3X1 U22506 ( .A(n24142), .B(n24645), .C(n22767), .Y(n21406) );
  AOI22X1 U22507 ( .A(n29408), .B(n26077), .C(n11949), .D(net96558), .Y(n33725) );
  MUX2X1 U22508 ( .B(n22714), .A(n29356), .S(n23467), .Y(n33723) );
  AOI21X1 U22509 ( .A(n29433), .B(n3147), .C(n33723), .Y(n33724) );
  AOI22X1 U22510 ( .A(n29399), .B(n26077), .C(n11948), .D(net96558), .Y(n33730) );
  MUX2X1 U22511 ( .B(n24296), .A(n29345), .S(n23467), .Y(n33728) );
  AOI21X1 U22512 ( .A(n29433), .B(n3146), .C(n33728), .Y(n33729) );
  AOI22X1 U22513 ( .A(n11947), .B(net96562), .C(n29407), .D(n33748), .Y(n33733) );
  AOI22X1 U22514 ( .A(n30519), .B(n29361), .C(n29414), .D(n26077), .Y(n33731)
         );
  NAND3X1 U22515 ( .A(n22645), .B(n24646), .C(n24834), .Y(n21401) );
  AOI22X1 U22516 ( .A(n30519), .B(n29351), .C(n29397), .D(n33748), .Y(n33736)
         );
  AOI22X1 U22517 ( .A(n11946), .B(net96562), .C(n29429), .D(n3144), .Y(n33734)
         );
  NAND3X1 U22518 ( .A(n24143), .B(n24647), .C(n22768), .Y(n21400) );
  AOI22X1 U22519 ( .A(n11945), .B(net96566), .C(n30519), .D(n29406), .Y(n33739) );
  AOI22X1 U22520 ( .A(n29361), .B(n26077), .C(n29414), .D(n33748), .Y(n33737)
         );
  NAND3X1 U22521 ( .A(n22646), .B(n24648), .C(n24835), .Y(n21398) );
  AOI22X1 U22522 ( .A(n29350), .B(n26077), .C(n30519), .D(n29396), .Y(n33742)
         );
  AOI22X1 U22523 ( .A(n11944), .B(net96562), .C(n29429), .D(n3142), .Y(n33740)
         );
  NAND3X1 U22524 ( .A(n24144), .B(n24649), .C(n22769), .Y(n21397) );
  AOI22X1 U22525 ( .A(n29408), .B(n33762), .C(n11943), .D(net96558), .Y(n33746) );
  MUX2X1 U22526 ( .B(n22715), .A(n29356), .S(n33748), .Y(n33744) );
  AOI21X1 U22527 ( .A(n29433), .B(n3141), .C(n33744), .Y(n33745) );
  AOI22X1 U22528 ( .A(n29399), .B(n33762), .C(n11942), .D(net96558), .Y(n33752) );
  MUX2X1 U22529 ( .B(n24297), .A(n29345), .S(n33748), .Y(n33750) );
  AOI21X1 U22530 ( .A(n29433), .B(n3140), .C(n33750), .Y(n33751) );
  AOI22X1 U22531 ( .A(n11941), .B(net96566), .C(n29407), .D(n23466), .Y(n33755) );
  AOI22X1 U22532 ( .A(n30514), .B(n29361), .C(n29414), .D(n33762), .Y(n33753)
         );
  NAND3X1 U22533 ( .A(n22647), .B(n24650), .C(n24836), .Y(n21392) );
  AOI22X1 U22534 ( .A(n30514), .B(n29351), .C(n29397), .D(n23466), .Y(n33758)
         );
  AOI22X1 U22535 ( .A(n11940), .B(net96566), .C(n29428), .D(n3138), .Y(n33756)
         );
  NAND3X1 U22536 ( .A(n24145), .B(n24651), .C(n22770), .Y(n21391) );
  AOI22X1 U22537 ( .A(n11939), .B(net96566), .C(n30514), .D(n29405), .Y(n33761) );
  AOI22X1 U22538 ( .A(n29359), .B(n33762), .C(n29414), .D(n23466), .Y(n33759)
         );
  NAND3X1 U22539 ( .A(n22648), .B(n24652), .C(n24837), .Y(n21389) );
  AOI22X1 U22540 ( .A(n29350), .B(n33762), .C(n30514), .D(n29396), .Y(n33765)
         );
  AOI22X1 U22541 ( .A(n11938), .B(net96566), .C(n29430), .D(n3136), .Y(n33763)
         );
  NAND3X1 U22542 ( .A(n24146), .B(n24653), .C(n22771), .Y(n21388) );
  AOI22X1 U22543 ( .A(n29409), .B(n33784), .C(n11937), .D(net96558), .Y(n33769) );
  MUX2X1 U22544 ( .B(n27046), .A(n29356), .S(n23466), .Y(n33767) );
  AOI21X1 U22545 ( .A(n29433), .B(n3135), .C(n33767), .Y(n33768) );
  AOI22X1 U22546 ( .A(n29399), .B(n33784), .C(n11936), .D(net96558), .Y(n33774) );
  MUX2X1 U22547 ( .B(n24298), .A(n29345), .S(n23466), .Y(n33772) );
  AOI21X1 U22548 ( .A(n29433), .B(n3134), .C(n33772), .Y(n33773) );
  AOI22X1 U22549 ( .A(n11935), .B(net96566), .C(n29408), .D(n25771), .Y(n33777) );
  AOI22X1 U22550 ( .A(n30509), .B(n29362), .C(n29414), .D(n33784), .Y(n33775)
         );
  NAND3X1 U22551 ( .A(n22649), .B(n24654), .C(n24838), .Y(n21383) );
  AOI22X1 U22552 ( .A(n30509), .B(n29351), .C(n29396), .D(n25771), .Y(n33780)
         );
  AOI22X1 U22553 ( .A(n11934), .B(net96564), .C(n29430), .D(n3132), .Y(n33778)
         );
  NAND3X1 U22554 ( .A(n24147), .B(n24655), .C(n22772), .Y(n21382) );
  AOI22X1 U22555 ( .A(n11933), .B(net96564), .C(n30509), .D(n29405), .Y(n33783) );
  AOI22X1 U22556 ( .A(n29361), .B(n33784), .C(n29414), .D(n25771), .Y(n33781)
         );
  NAND3X1 U22557 ( .A(n22650), .B(n24656), .C(n24839), .Y(n21380) );
  AOI22X1 U22558 ( .A(n29350), .B(n33784), .C(n30509), .D(n29396), .Y(n33787)
         );
  AOI22X1 U22559 ( .A(n11932), .B(net96564), .C(n29430), .D(n3130), .Y(n33785)
         );
  NAND3X1 U22560 ( .A(n24148), .B(n24657), .C(n22773), .Y(n21379) );
  AOI22X1 U22561 ( .A(n29409), .B(n33806), .C(n11931), .D(net96558), .Y(n33791) );
  MUX2X1 U22562 ( .B(n27045), .A(n29356), .S(n25771), .Y(n33789) );
  AOI21X1 U22563 ( .A(n29433), .B(n3129), .C(n33789), .Y(n33790) );
  AOI22X1 U22564 ( .A(n29399), .B(n33806), .C(n11930), .D(net96558), .Y(n33796) );
  MUX2X1 U22565 ( .B(n26899), .A(n29345), .S(n25771), .Y(n33794) );
  AOI21X1 U22566 ( .A(n29433), .B(n3128), .C(n33794), .Y(n33795) );
  AOI22X1 U22567 ( .A(n30504), .B(n29362), .C(n29407), .D(n33815), .Y(n33799)
         );
  AOI22X1 U22568 ( .A(n11929), .B(net96564), .C(n29430), .D(n3127), .Y(n33797)
         );
  NAND3X1 U22569 ( .A(n24149), .B(n24658), .C(n22774), .Y(n21374) );
  AOI22X1 U22570 ( .A(n30504), .B(n29351), .C(n29396), .D(n33815), .Y(n33802)
         );
  AOI22X1 U22571 ( .A(n11928), .B(net96564), .C(n29430), .D(n3126), .Y(n33800)
         );
  NAND3X1 U22572 ( .A(n24150), .B(n24659), .C(n22775), .Y(n21373) );
  AOI22X1 U22573 ( .A(n29361), .B(n33806), .C(n30504), .D(n29405), .Y(n33805)
         );
  AOI22X1 U22574 ( .A(n11927), .B(net96564), .C(n29430), .D(n3125), .Y(n33803)
         );
  NAND3X1 U22575 ( .A(n24151), .B(n24660), .C(n22776), .Y(n21371) );
  AOI22X1 U22576 ( .A(n29350), .B(n33806), .C(n30504), .D(n29397), .Y(n33809)
         );
  AOI22X1 U22577 ( .A(n11926), .B(net96568), .C(n29431), .D(n26071), .Y(n33807) );
  NAND3X1 U22578 ( .A(n24152), .B(n24661), .C(n22777), .Y(n21370) );
  AOI22X1 U22579 ( .A(n29409), .B(n33829), .C(n11925), .D(net96558), .Y(n33813) );
  MUX2X1 U22580 ( .B(n22716), .A(n29356), .S(n33815), .Y(n33811) );
  AOI21X1 U22581 ( .A(n29433), .B(n3123), .C(n33811), .Y(n33812) );
  AOI22X1 U22582 ( .A(n29400), .B(n25675), .C(n11924), .D(net96558), .Y(n33819) );
  MUX2X1 U22583 ( .B(n24299), .A(n29345), .S(n33815), .Y(n33817) );
  AOI21X1 U22584 ( .A(n29432), .B(n3122), .C(n33817), .Y(n33818) );
  AOI22X1 U22585 ( .A(n23292), .B(n29362), .C(n29406), .D(n25830), .Y(n33822)
         );
  AOI22X1 U22586 ( .A(n11923), .B(net96568), .C(n29430), .D(n3121), .Y(n33820)
         );
  NAND3X1 U22587 ( .A(n24153), .B(n24662), .C(n22778), .Y(n21365) );
  AOI22X1 U22588 ( .A(n23292), .B(n29351), .C(n29396), .D(n25830), .Y(n33825)
         );
  AOI22X1 U22589 ( .A(n11922), .B(net96568), .C(n29430), .D(n3120), .Y(n33823)
         );
  NAND3X1 U22590 ( .A(n24154), .B(n24663), .C(n22779), .Y(n21364) );
  AOI22X1 U22591 ( .A(n29360), .B(n25675), .C(n23292), .D(n29405), .Y(n33828)
         );
  AOI22X1 U22592 ( .A(n11921), .B(net96568), .C(n29430), .D(n3119), .Y(n33826)
         );
  NAND3X1 U22593 ( .A(n24155), .B(n24664), .C(n22780), .Y(n21362) );
  AOI22X1 U22594 ( .A(n29350), .B(n33829), .C(n23292), .D(n29396), .Y(n33832)
         );
  AOI22X1 U22595 ( .A(n11920), .B(net96568), .C(n29429), .D(n3118), .Y(n33830)
         );
  NAND3X1 U22596 ( .A(n24156), .B(n24665), .C(n22781), .Y(n21361) );
  AOI22X1 U22597 ( .A(n29408), .B(n33852), .C(n11919), .D(net96558), .Y(n33836) );
  MUX2X1 U22598 ( .B(n26900), .A(n29356), .S(n25830), .Y(n33834) );
  AOI21X1 U22599 ( .A(n29432), .B(n3117), .C(n33834), .Y(n33835) );
  AOI22X1 U22600 ( .A(n29400), .B(n33852), .C(n11918), .D(net96558), .Y(n33841) );
  MUX2X1 U22601 ( .B(n24300), .A(n29345), .S(n25830), .Y(n33839) );
  AOI21X1 U22602 ( .A(n29432), .B(n3116), .C(n33839), .Y(n33840) );
  AOI22X1 U22603 ( .A(n30495), .B(n29362), .C(n29406), .D(n33861), .Y(n33845)
         );
  AOI22X1 U22604 ( .A(n11917), .B(net96568), .C(n29429), .D(n3115), .Y(n33843)
         );
  NAND3X1 U22605 ( .A(n24157), .B(n24666), .C(n22782), .Y(n21356) );
  AOI22X1 U22606 ( .A(n30495), .B(n29351), .C(n29397), .D(n33861), .Y(n33848)
         );
  AOI22X1 U22607 ( .A(n11916), .B(net96568), .C(n29430), .D(n3114), .Y(n33846)
         );
  NAND3X1 U22608 ( .A(n24158), .B(n24667), .C(n22783), .Y(n21355) );
  AOI22X1 U22609 ( .A(n29361), .B(n33852), .C(n30495), .D(n29405), .Y(n33851)
         );
  AOI22X1 U22610 ( .A(n11915), .B(net96566), .C(n29430), .D(n3113), .Y(n33849)
         );
  NAND3X1 U22611 ( .A(n24159), .B(n24668), .C(n22784), .Y(n21353) );
  AOI22X1 U22612 ( .A(n29350), .B(n33852), .C(n30495), .D(n29396), .Y(n33855)
         );
  AOI22X1 U22613 ( .A(n11914), .B(net96566), .C(n29430), .D(n3112), .Y(n33853)
         );
  NAND3X1 U22614 ( .A(n24160), .B(n24669), .C(n22785), .Y(n21352) );
  AOI22X1 U22615 ( .A(n29409), .B(n33875), .C(n11913), .D(net96558), .Y(n33859) );
  MUX2X1 U22616 ( .B(n26965), .A(n29356), .S(n33861), .Y(n33857) );
  AOI21X1 U22617 ( .A(n29432), .B(n3111), .C(n33857), .Y(n33858) );
  AOI22X1 U22618 ( .A(n29400), .B(n33875), .C(n11912), .D(net96558), .Y(n33865) );
  MUX2X1 U22619 ( .B(n26898), .A(n29345), .S(n33861), .Y(n33863) );
  AOI21X1 U22620 ( .A(n29432), .B(n3110), .C(n33863), .Y(n33864) );
  AOI22X1 U22621 ( .A(n23287), .B(n29361), .C(n29407), .D(n33884), .Y(n33868)
         );
  AOI22X1 U22622 ( .A(n11911), .B(net96566), .C(n29430), .D(n25751), .Y(n33866) );
  NAND3X1 U22623 ( .A(n24161), .B(n24670), .C(n22786), .Y(n21347) );
  AOI22X1 U22624 ( .A(n23287), .B(n29351), .C(n29396), .D(n33884), .Y(n33871)
         );
  AOI22X1 U22625 ( .A(n11910), .B(net96566), .C(n29429), .D(n3108), .Y(n33869)
         );
  NAND3X1 U22626 ( .A(n24162), .B(n24671), .C(n22787), .Y(n21346) );
  AOI22X1 U22627 ( .A(n29360), .B(n33875), .C(n23287), .D(n29405), .Y(n33874)
         );
  AOI22X1 U22628 ( .A(n11909), .B(net96566), .C(n29429), .D(n3107), .Y(n33872)
         );
  NAND3X1 U22629 ( .A(n24163), .B(n24672), .C(n22788), .Y(n21344) );
  AOI22X1 U22630 ( .A(n29350), .B(n33875), .C(n23287), .D(n29400), .Y(n33878)
         );
  AOI22X1 U22631 ( .A(n11908), .B(net96566), .C(n29429), .D(n3106), .Y(n33876)
         );
  NAND3X1 U22632 ( .A(n24164), .B(n24673), .C(n22789), .Y(n21343) );
  AOI22X1 U22633 ( .A(n29409), .B(n33900), .C(n11907), .D(net96558), .Y(n33882) );
  MUX2X1 U22634 ( .B(n22717), .A(n29356), .S(n33884), .Y(n33880) );
  AOI21X1 U22635 ( .A(n29432), .B(n3105), .C(n33880), .Y(n33881) );
  AOI22X1 U22636 ( .A(n29399), .B(n33900), .C(n11906), .D(net96558), .Y(n33889) );
  MUX2X1 U22637 ( .B(n22718), .A(n29345), .S(n33884), .Y(n33887) );
  AOI21X1 U22638 ( .A(n29432), .B(n3104), .C(n33887), .Y(n33888) );
  AOI22X1 U22639 ( .A(n33890), .B(n29361), .C(n29407), .D(n33908), .Y(n33893)
         );
  AOI22X1 U22640 ( .A(n11905), .B(net96566), .C(n29429), .D(n3103), .Y(n33891)
         );
  NAND3X1 U22641 ( .A(n24165), .B(n24674), .C(n22790), .Y(n21338) );
  AOI22X1 U22642 ( .A(n33890), .B(n29351), .C(n29397), .D(n33908), .Y(n33896)
         );
  AOI22X1 U22643 ( .A(n11904), .B(net96570), .C(n29429), .D(n3102), .Y(n33894)
         );
  NAND3X1 U22644 ( .A(n24166), .B(n24675), .C(n22791), .Y(n21337) );
  AOI22X1 U22645 ( .A(n29360), .B(n33900), .C(n33890), .D(n29405), .Y(n33899)
         );
  AOI22X1 U22646 ( .A(n11903), .B(net96570), .C(data_in[5]), .D(n29424), .Y(
        n33897) );
  NAND3X1 U22647 ( .A(n24167), .B(n24676), .C(n22792), .Y(n21335) );
  AOI22X1 U22648 ( .A(n29350), .B(n33900), .C(n33890), .D(n29399), .Y(n33903)
         );
  AOI22X1 U22649 ( .A(n11902), .B(net96568), .C(data_in[4]), .D(n29424), .Y(
        n33901) );
  NAND3X1 U22650 ( .A(n24168), .B(n24677), .C(n22793), .Y(n21334) );
  AOI22X1 U22651 ( .A(n29360), .B(n33908), .C(n23275), .D(n29405), .Y(n33907)
         );
  AOI22X1 U22652 ( .A(net96570), .B(n11901), .C(data_in[3]), .D(n29424), .Y(
        n33905) );
  NAND3X1 U22653 ( .A(n24169), .B(n24678), .C(n20959), .Y(n21332) );
  AOI22X1 U22654 ( .A(n29350), .B(n33908), .C(n23275), .D(n29398), .Y(n33911)
         );
  AOI22X1 U22655 ( .A(n11900), .B(net96568), .C(data_in[2]), .D(n29424), .Y(
        n33909) );
  NAND3X1 U22656 ( .A(n24170), .B(n24679), .C(n24841), .Y(n21331) );
  AOI22X1 U22657 ( .A(n12024), .B(net96568), .C(n30577), .D(n29348), .Y(n33915) );
  AOI22X1 U22658 ( .A(n29399), .B(n20856), .C(n29429), .D(n3222), .Y(n33913)
         );
  NAND3X1 U22659 ( .A(n24842), .B(n24680), .C(n22651), .Y(n21518) );
  NAND2X1 U22660 ( .A(n30656), .B(n33992), .Y(n33916) );
  NAND3X1 U22661 ( .A(n19663), .B(n33917), .C(n33919), .Y(n34179) );
  NAND3X1 U22662 ( .A(n33917), .B(n33920), .C(n19664), .Y(n34178) );
  NAND3X1 U22663 ( .A(n33917), .B(n19664), .C(n19663), .Y(n33918) );
  NAND3X1 U22664 ( .A(n19662), .B(n33920), .C(n33919), .Y(n34213) );
  MUX2X1 U22665 ( .B(n25615), .A(n20994), .S(n27296), .Y(n33921) );
  OAI21X1 U22666 ( .A(n21044), .B(n26076), .C(n33921), .Y(n33922) );
  AOI22X1 U22667 ( .A(n23280), .B(n33922), .C(n27309), .D(n27912), .Y(n33925)
         );
  AOI22X1 U22668 ( .A(n27267), .B(net105798), .C(n29352), .D(n23611), .Y(
        n33924) );
  MUX2X1 U22669 ( .B(n22719), .A(n21044), .S(alt5_net95664), .Y(n33927) );
  AOI22X1 U22670 ( .A(n27267), .B(net110825), .C(n29352), .D(n21007), .Y(
        n33929) );
  NAND3X1 U22671 ( .A(wS), .B(n34504), .C(n34497), .Y(n33931) );
  NAND2X1 U22672 ( .A(n15201), .B(n33931), .Y(n22326) );
  NAND2X1 U22673 ( .A(n25338), .B(n33992), .Y(n33932) );
  OAI21X1 U22674 ( .A(net151875), .B(net90055), .C(n23209), .Y(net90054) );
  AOI22X1 U22675 ( .A(n4218), .B(net147500), .C(n3304), .D(net110809), .Y(
        n33936) );
  AOI22X1 U22676 ( .A(n4217), .B(net147499), .C(n3303), .D(net117217), .Y(
        n33938) );
  AOI22X1 U22677 ( .A(n4216), .B(net147496), .C(n3302), .D(net107078), .Y(
        n33940) );
  AOI22X1 U22678 ( .A(n4215), .B(net147501), .C(n3301), .D(net107094), .Y(
        n33942) );
  AOI22X1 U22679 ( .A(n4214), .B(net147504), .C(n3300), .D(net117217), .Y(
        n33944) );
  AOI22X1 U22680 ( .A(n4213), .B(net147507), .C(n3299), .D(net107090), .Y(
        n33946) );
  AOI22X1 U22681 ( .A(n4212), .B(net147498), .C(n3298), .D(n20851), .Y(n33948)
         );
  AOI22X1 U22682 ( .A(n4211), .B(net147499), .C(n3297), .D(net107082), .Y(
        n33950) );
  AOI22X1 U22683 ( .A(n4210), .B(net147497), .C(n3296), .D(net151840), .Y(
        n33952) );
  AOI22X1 U22684 ( .A(n4209), .B(net147502), .C(n3295), .D(net107094), .Y(
        n33954) );
  AOI22X1 U22685 ( .A(n4207), .B(net147501), .C(n3293), .D(net107061), .Y(
        n33956) );
  AOI22X1 U22686 ( .A(n4206), .B(net147498), .C(n3292), .D(n20854), .Y(n33958)
         );
  AOI22X1 U22687 ( .A(n4205), .B(net147502), .C(n3291), .D(net107061), .Y(
        n33960) );
  AOI22X1 U22688 ( .A(n4204), .B(net147499), .C(n3290), .D(net150376), .Y(
        n33962) );
  AOI22X1 U22689 ( .A(n4203), .B(net147505), .C(n3289), .D(net107090), .Y(
        n33964) );
  AOI22X1 U22690 ( .A(n4202), .B(net147502), .C(n3288), .D(net107061), .Y(
        n33966) );
  AOI22X1 U22691 ( .A(n4201), .B(net147505), .C(n3287), .D(net151649), .Y(
        n33968) );
  AOI22X1 U22692 ( .A(n4200), .B(net151738), .C(n3286), .D(net151814), .Y(
        n33970) );
  AOI22X1 U22693 ( .A(n4198), .B(net147501), .C(n3284), .D(n20854), .Y(n33973)
         );
  AOI22X1 U22694 ( .A(n4197), .B(net147506), .C(n3283), .D(net107090), .Y(
        n33975) );
  AOI22X1 U22695 ( .A(n4196), .B(net151738), .C(n3282), .D(net150376), .Y(
        n33977) );
  AOI22X1 U22696 ( .A(n4195), .B(net147497), .C(n3281), .D(net151814), .Y(
        n33979) );
  AOI22X1 U22697 ( .A(n4194), .B(net151751), .C(n3280), .D(net150376), .Y(
        n33981) );
  AOI22X1 U22698 ( .A(n4193), .B(net147507), .C(n3279), .D(net107088), .Y(
        n33983) );
  AOI22X1 U22699 ( .A(n4192), .B(net147504), .C(n3278), .D(net107082), .Y(
        n33985) );
  AOI22X1 U22700 ( .A(n4191), .B(net151751), .C(n3277), .D(net107063), .Y(
        n33987) );
  AOI22X1 U22701 ( .A(n4219), .B(net147507), .C(n3305), .D(net151649), .Y(
        n33989) );
  AOI22X1 U22702 ( .A(n4190), .B(net151738), .C(n3276), .D(net107088), .Y(
        n33991) );
  NAND3X1 U22703 ( .A(n21204), .B(net114546), .C(n33992), .Y(n33994) );
  NAND2X1 U22704 ( .A(n15201), .B(n15204), .Y(n22324) );
  AND2X2 U22705 ( .A(n9127), .B(n29380), .Y(n21784) );
  AND2X2 U22706 ( .A(n9128), .B(n29381), .Y(n21785) );
  AND2X2 U22707 ( .A(n9129), .B(n29381), .Y(n21786) );
  AND2X2 U22708 ( .A(n9131), .B(n29381), .Y(n21788) );
  AND2X2 U22709 ( .A(n9139), .B(n29381), .Y(n21796) );
  AND2X2 U22710 ( .A(n9143), .B(n29380), .Y(n21800) );
  AND2X2 U22711 ( .A(n9145), .B(n29381), .Y(n21803) );
  AND2X2 U22712 ( .A(n9147), .B(n29381), .Y(n21805) );
  AND2X2 U22713 ( .A(n9148), .B(n29381), .Y(n21806) );
  AND2X2 U22714 ( .A(n9149), .B(n29381), .Y(n21807) );
  AND2X2 U22715 ( .A(n9151), .B(n29381), .Y(n21809) );
  AND2X2 U22716 ( .A(n9152), .B(n29381), .Y(n21810) );
  AND2X2 U22717 ( .A(n9153), .B(n29381), .Y(n21811) );
  AND2X2 U22718 ( .A(n9154), .B(n29381), .Y(n21812) );
  AND2X2 U22719 ( .A(n9155), .B(n29381), .Y(n21813) );
  NAND3X1 U22720 ( .A(n34171), .B(n25778), .C(n34170), .Y(n34176) );
  NAND3X1 U22721 ( .A(n13802), .B(n25686), .C(n24873), .Y(n34175) );
  OAI21X1 U22722 ( .A(n22686), .B(n24687), .C(n24973), .Y(n21323) );
  AOI22X1 U22723 ( .A(n20999), .B(n27186), .C(n34196), .D(n27318), .Y(n34181)
         );
  MUX2X1 U22724 ( .B(n34199), .A(n34198), .S(n27297), .Y(n34180) );
  AOI22X1 U22725 ( .A(n23280), .B(n22724), .C(n27309), .D(n25688), .Y(n34184)
         );
  AOI22X1 U22726 ( .A(n27267), .B(net104479), .C(n30078), .D(n21217), .Y(
        n34183) );
  AOI22X1 U22727 ( .A(n29185), .B(n34211), .C(n25615), .D(n26164), .Y(n34186)
         );
  AOI22X1 U22728 ( .A(n23280), .B(n22723), .C(n27309), .D(n27915), .Y(n34191)
         );
  AOI22X1 U22729 ( .A(n27267), .B(net149862), .C(n30078), .D(n23441), .Y(
        n34190) );
  AOI22X1 U22730 ( .A(n27241), .B(n29351), .C(n34192), .D(n29397), .Y(n34195)
         );
  AOI22X1 U22731 ( .A(n11898), .B(net96568), .C(data_in[0]), .D(n29424), .Y(
        n34193) );
  NAND3X1 U22732 ( .A(n22652), .B(n24681), .C(n24844), .Y(n21328) );
  AOI22X1 U22733 ( .A(n20999), .B(n34197), .C(n20994), .D(n27317), .Y(n34201)
         );
  AOI22X1 U22734 ( .A(n34199), .B(n27320), .C(n34198), .D(n27321), .Y(n34200)
         );
  AOI22X1 U22735 ( .A(n23280), .B(n24316), .C(n27309), .D(n20969), .Y(n34205)
         );
  AOI22X1 U22736 ( .A(n27267), .B(net124030), .C(n29352), .D(n26339), .Y(
        n34204) );
  AOI22X1 U22737 ( .A(n27241), .B(n29362), .C(n34192), .D(n29405), .Y(n34208)
         );
  AOI22X1 U22738 ( .A(n11899), .B(net96568), .C(data_in[1]), .D(n29424), .Y(
        n34206) );
  NAND3X1 U22739 ( .A(n23609), .B(n24682), .C(n24846), .Y(n21329) );
  AOI22X1 U22740 ( .A(n34211), .B(n34210), .C(n25615), .D(n25731), .Y(n34212)
         );
  OAI21X1 U22741 ( .A(net89744), .B(n21029), .C(n21924), .Y(n34214) );
  AOI22X1 U22742 ( .A(n23280), .B(n34214), .C(n27309), .D(n25649), .Y(n34217)
         );
  AOI22X1 U22743 ( .A(n27267), .B(n28220), .C(n30078), .D(n21183), .Y(n34216)
         );
  MUX2X1 U22744 ( .B(n22720), .A(n29356), .S(n34342), .Y(n34221) );
  AOI21X1 U22745 ( .A(n29408), .B(n34222), .C(n34221), .Y(n34223) );
  OAI21X1 U22746 ( .A(n34225), .B(n29212), .C(n23883), .Y(n34226) );
  AOI22X1 U22747 ( .A(n34228), .B(n34227), .C(n34228), .D(net96596), .Y(n34460) );
  NAND3X1 U22748 ( .A(n21104), .B(n34279), .C(n34230), .Y(n34437) );
  AOI21X1 U22749 ( .A(T[4]), .B(n34355), .C(n25725), .Y(n34236) );
  OAI21X1 U22750 ( .A(n34235), .B(n34351), .C(n23000), .Y(n34244) );
  OAI21X1 U22751 ( .A(n34243), .B(n24689), .C(n34242), .Y(n34237) );
  OAI21X1 U22752 ( .A(n22973), .B(n34305), .C(n26057), .Y(n34240) );
  OAI21X1 U22753 ( .A(n25759), .B(n34264), .C(n34240), .Y(n34262) );
  OAI21X1 U22754 ( .A(n34243), .B(n25326), .C(n25222), .Y(n34250) );
  AOI21X1 U22755 ( .A(n25223), .B(n25126), .C(n22274), .Y(n34247) );
  AOI21X1 U22756 ( .A(n25689), .B(n21523), .C(n34261), .Y(n34253) );
  NAND3X1 U22757 ( .A(n23187), .B(n23000), .C(n34250), .Y(n34256) );
  XNOR2X1 U22758 ( .A(n23105), .B(n25160), .Y(n34254) );
  XNOR2X1 U22759 ( .A(n34254), .B(n25169), .Y(n34278) );
  NAND3X1 U22760 ( .A(n21523), .B(n25317), .C(n25689), .Y(n34258) );
  OAI21X1 U22761 ( .A(n34261), .B(n25317), .C(n21986), .Y(n34276) );
  OAI21X1 U22762 ( .A(n25004), .B(n34260), .C(n34315), .Y(n34275) );
  AOI21X1 U22763 ( .A(n34270), .B(n34407), .C(n34326), .Y(n34268) );
  OAI21X1 U22764 ( .A(n23071), .B(n25446), .C(n22973), .Y(n34267) );
  OAI21X1 U22765 ( .A(n25766), .B(n20963), .C(n21993), .Y(n34271) );
  AOI22X1 U22766 ( .A(n25862), .B(n34273), .C(n21524), .D(n34271), .Y(n34274)
         );
  OAI21X1 U22767 ( .A(n34276), .B(n34275), .C(n21925), .Y(n34277) );
  OAI21X1 U22768 ( .A(n26055), .B(n34278), .C(n34277), .Y(n34281) );
  AOI22X1 U22769 ( .A(n29387), .B(n34342), .C(n29351), .D(n23457), .Y(n34285)
         );
  AOI22X1 U22770 ( .A(n29432), .B(n3274), .C(n29397), .D(n23424), .Y(n34284)
         );
  AND2X2 U22771 ( .A(n23587), .B(n23738), .Y(n34287) );
  AOI22X1 U22772 ( .A(n34287), .B(n34286), .C(n34287), .D(net96596), .Y(n34493) );
  AOI22X1 U22773 ( .A(n4220), .B(net147496), .C(n3306), .D(net107061), .Y(
        n34289) );
  OAI21X1 U22774 ( .A(n25688), .B(n22733), .C(n34441), .Y(n34290) );
  OAI21X1 U22775 ( .A(n34351), .B(n34291), .C(n23001), .Y(n34295) );
  OAI21X1 U22776 ( .A(n25630), .B(n25324), .C(n21988), .Y(n34310) );
  AOI21X1 U22777 ( .A(n25834), .B(n22679), .C(n22278), .Y(n34299) );
  AOI21X1 U22778 ( .A(T[4]), .B(n25688), .C(n34302), .Y(n34297) );
  OAI21X1 U22779 ( .A(n22687), .B(n26046), .C(n25668), .Y(n34298) );
  MUX2X1 U22780 ( .B(n22721), .A(n24320), .S(n26065), .Y(n34301) );
  INVX2 U22781 ( .A(n34301), .Y(n34322) );
  MUX2X1 U22782 ( .B(n25324), .A(n34302), .S(n26049), .Y(n34304) );
  OAI21X1 U22783 ( .A(n34305), .B(n25435), .C(n25850), .Y(n34306) );
  OAI21X1 U22784 ( .A(n25759), .B(n34307), .C(n34306), .Y(n34321) );
  NAND3X1 U22785 ( .A(n23001), .B(n26064), .C(n34310), .Y(n34316) );
  OAI21X1 U22786 ( .A(n26055), .B(n34314), .C(n25580), .Y(n34340) );
  AOI21X1 U22787 ( .A(n34320), .B(n25225), .C(n34434), .Y(n34337) );
  AOI22X1 U22788 ( .A(n34318), .B(n27074), .C(n34319), .D(n25225), .Y(n34336)
         );
  FAX1 U22789 ( .A(n34323), .B(n34322), .C(n34321), .YC(), .YS(n34334) );
  FAX1 U22790 ( .A(n25759), .B(n25436), .C(n25850), .YC(), .YS(n34330) );
  OAI21X1 U22791 ( .A(n23073), .B(n25446), .C(n25435), .Y(n34328) );
  OAI21X1 U22792 ( .A(n25766), .B(n34330), .C(n34329), .Y(n34331) );
  OAI21X1 U22793 ( .A(n25862), .B(n34332), .C(n34331), .Y(n34333) );
  OAI21X1 U22794 ( .A(n34417), .B(n34334), .C(n34333), .Y(n34335) );
  AOI21X1 U22795 ( .A(n24261), .B(n24245), .C(n34335), .Y(n34339) );
  AOI22X1 U22796 ( .A(n29407), .B(n23424), .C(n29429), .D(n3275), .Y(n34345)
         );
  AOI22X1 U22797 ( .A(n29360), .B(n23457), .C(n29414), .D(n34342), .Y(n34344)
         );
  AOI22X1 U22798 ( .A(n27283), .B(n34346), .C(n27283), .D(net96596), .Y(n34494) );
  AOI22X1 U22799 ( .A(n4221), .B(net147505), .C(n3307), .D(net107088), .Y(
        n34348) );
  AND2X2 U22800 ( .A(n9157), .B(n29381), .Y(n21815) );
  NOR3X1 U22801 ( .A(n34443), .B(n23274), .C(n22938), .Y(n34350) );
  OAI21X1 U22802 ( .A(n25838), .B(n34351), .C(n27158), .Y(n34367) );
  XOR2X1 U22803 ( .A(n34353), .B(n25636), .Y(n34361) );
  NAND3X1 U22804 ( .A(n26054), .B(n34354), .C(T[3]), .Y(n34403) );
  AOI21X1 U22805 ( .A(n34358), .B(n22993), .C(n25844), .Y(n34359) );
  OAI21X1 U22806 ( .A(n34362), .B(n34361), .C(n34360), .Y(n34402) );
  NAND3X1 U22807 ( .A(n26058), .B(n22993), .C(n24874), .Y(n34370) );
  AOI21X1 U22808 ( .A(n27295), .B(n34390), .C(n34365), .Y(n34368) );
  OAI21X1 U22809 ( .A(n34367), .B(n24691), .C(n27158), .Y(n34369) );
  MUX2X1 U22810 ( .B(n24301), .A(n24321), .S(n25667), .Y(n34426) );
  XOR2X1 U22811 ( .A(n20967), .B(n25661), .Y(n34374) );
  OAI21X1 U22812 ( .A(n25863), .B(n25405), .C(n23888), .Y(n34422) );
  AOI21X1 U22813 ( .A(n34378), .B(n20967), .C(n21399), .Y(n34377) );
  OAI21X1 U22814 ( .A(n34378), .B(n21226), .C(n21987), .Y(n34382) );
  XOR2X1 U22815 ( .A(n34422), .B(n20970), .Y(n34389) );
  NAND3X1 U22816 ( .A(n22672), .B(n34391), .C(n25851), .Y(n34388) );
  AOI21X1 U22817 ( .A(T[1]), .B(n25661), .C(n25664), .Y(n34384) );
  OAI21X1 U22818 ( .A(n25863), .B(n25133), .C(n34383), .Y(n34387) );
  MUX2X1 U22819 ( .B(n34389), .A(n24322), .S(n25681), .Y(n34425) );
  OAI21X1 U22820 ( .A(n34390), .B(n34358), .C(n21525), .Y(n34411) );
  XOR2X1 U22821 ( .A(n25752), .B(n25322), .Y(n34405) );
  XOR2X1 U22822 ( .A(n25417), .B(n21228), .Y(n34397) );
  OAI21X1 U22823 ( .A(n25780), .B(n34411), .C(n25734), .Y(n34398) );
  OAI21X1 U22824 ( .A(n34400), .B(n34405), .C(n34398), .Y(n34423) );
  FAX1 U22825 ( .A(n25748), .B(n34399), .C(n25750), .YC(), .YS(n34418) );
  FAX1 U22826 ( .A(n34404), .B(n21124), .C(n34400), .YC(), .YS(n34415) );
  NAND3X1 U22827 ( .A(n34401), .B(n25416), .C(n34402), .Y(n34412) );
  NAND3X1 U22828 ( .A(n25858), .B(n34405), .C(n34406), .Y(n34409) );
  NAND3X1 U22829 ( .A(n25858), .B(n25780), .C(n25860), .Y(n34408) );
  AOI21X1 U22830 ( .A(n34415), .B(n34414), .C(n34413), .Y(n34416) );
  AOI21X1 U22831 ( .A(n34417), .B(n34418), .C(n22146), .Y(n34419) );
  NAND3X1 U22832 ( .A(n22974), .B(n26059), .C(n34432), .Y(n34430) );
  AOI21X1 U22833 ( .A(n34431), .B(n23277), .C(n34434), .Y(n34428) );
  NAND3X1 U22834 ( .A(n24237), .B(n24683), .C(n24856), .Y(n34439) );
  AOI21X1 U22835 ( .A(n24265), .B(n34440), .C(n34438), .Y(n11043) );
  INVX2 U22840 ( .A(n2219), .Y(n14373) );
endmodule


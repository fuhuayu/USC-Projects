module lifo (
	push, 
	pop, 
	reset, 
	clk, 
	din, 
	empty, 
	full, 
	dout);
   input push;
   input pop;
   input reset;
   input clk;
   input [15:0] din;
   output empty;
   output full;
   output [15:0] dout;

   // Internal wires
   wire FE_PHN82_mem_16_;
   wire FE_PHN81_mem_47_;
   wire FE_PHN80_mem_71_;
   wire FE_PHN79_mem_119_;
   wire FE_PHN78_mem_27_;
   wire FE_PHN77_mem_31_;
   wire FE_PHN76_mem_19_;
   wire FE_PHN75_mem_20_;
   wire FE_PHN74_n247;
   wire FE_PHN73_mem_28_;
   wire FE_PHN72_mem_23_;
   wire FE_PHN71_mem_30_;
   wire FE_PHN70_mem_29_;
   wire FE_PHN69_mem_16_;
   wire FE_PHN68_mem_26_;
   wire FE_PHN67_n726;
   wire FE_PHN66_n686;
   wire FE_PHN65_FE_OFCN5_n231;
   wire FE_PHN64_FE_OFCN14_n222;
   wire FE_PHN63_FE_OFCN12_n224;
   wire FE_PHN62_FE_OFCN15_n221;
   wire FE_PHN61_FE_OFCN10_n226;
   wire FE_PHN60_FE_OFCN7_n229;
   wire FE_PHN59_FE_OFCN11_n225;
   wire FE_PHN58_FE_OFCN13_n223;
   wire FE_PHN57_FE_OFCN8_n228;
   wire FE_PHN56_FE_OFCN5_n231;
   wire FE_PHN55_FE_OFCN16_n219;
   wire FE_PHN54_FE_OFCN14_n222;
   wire FE_PHN53_FE_OFCN6_n230;
   wire FE_PHN52_FE_OFCN2_n234;
   wire FE_PHN51_FE_OFCN4_n232;
   wire FE_PHN50_FE_OFCN3_n233;
   wire FE_PHN49_FE_OFCN1_n235;
   wire FE_PHN48_FE_OFCN9_n227;
   wire FE_PSN47_n686;
   wire FE_PSN46_n34;
   wire FE_PSN45_full;
   wire FE_PSN44_n36;
   wire FE_PSN43_n36;
   wire FE_PSN42_FE_OFCN26_n105;
   wire FE_PSN41_FE_OFCN28_n123;
   wire FE_PSN40_n708;
   wire FE_PSN39_FE_OFCN28_n123;
   wire FE_PSN38_FE_OFCN29_n55;
   wire FE_PSN37_n55;
   wire FE_PSN36_FE_OFCN28_n123;
   wire FE_OFCN29_n55;
   wire FE_OFCN28_n123;
   wire FE_OFCN26_n105;
   wire FE_OFCN20_n199;
   wire FE_OFCN19_n239;
   wire FE_OFCN18_n245;
   wire FE_OFCN17_n241;
   wire FE_OFCN16_n219;
   wire FE_OFCN15_n221;
   wire FE_OFCN14_n222;
   wire FE_OFCN13_n223;
   wire FE_OFCN12_n224;
   wire FE_OFCN11_n225;
   wire FE_OFCN10_n226;
   wire FE_OFCN9_n227;
   wire FE_OFCN8_n228;
   wire FE_OFCN7_n229;
   wire FE_OFCN6_n230;
   wire FE_OFCN5_n231;
   wire FE_OFCN4_n232;
   wire FE_OFCN3_n233;
   wire FE_OFCN2_n234;
   wire FE_OFCN1_n235;
   wire clk__L2_N3;
   wire clk__L2_N2;
   wire clk__L2_N1;
   wire clk__L2_N0;
   wire clk__L1_N0;
   wire n34;
   wire n35;
   wire n36;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire [127:0] mem;

   BUFX2 FE_PHC82_mem_16_ (.Y(FE_PHN82_mem_16_), 
	.A(FE_PHN69_mem_16_));
   CLKBUF3 FE_PHC81_mem_47_ (.Y(FE_PHN81_mem_47_), 
	.A(mem[47]));
   CLKBUF2 FE_PHC80_mem_71_ (.Y(FE_PHN80_mem_71_), 
	.A(mem[71]));
   CLKBUF2 FE_PHC79_mem_119_ (.Y(FE_PHN79_mem_119_), 
	.A(mem[119]));
   CLKBUF2 FE_PHC78_mem_27_ (.Y(FE_PHN78_mem_27_), 
	.A(mem[27]));
   CLKBUF2 FE_PHC77_mem_31_ (.Y(FE_PHN77_mem_31_), 
	.A(mem[31]));
   CLKBUF2 FE_PHC76_mem_19_ (.Y(FE_PHN76_mem_19_), 
	.A(mem[19]));
   CLKBUF2 FE_PHC75_mem_20_ (.Y(FE_PHN75_mem_20_), 
	.A(mem[20]));
   BUFX2 FE_PHC74_n247 (.Y(FE_PHN74_n247), 
	.A(n247));
   CLKBUF2 FE_PHC73_mem_28_ (.Y(FE_PHN73_mem_28_), 
	.A(mem[28]));
   BUFX2 FE_PHC72_mem_23_ (.Y(FE_PHN72_mem_23_), 
	.A(mem[23]));
   BUFX2 FE_PHC71_mem_30_ (.Y(FE_PHN71_mem_30_), 
	.A(mem[30]));
   BUFX2 FE_PHC70_mem_29_ (.Y(FE_PHN70_mem_29_), 
	.A(mem[29]));
   BUFX2 FE_PHC69_mem_16_ (.Y(FE_PHN69_mem_16_), 
	.A(mem[16]));
   BUFX2 FE_PHC68_mem_26_ (.Y(FE_PHN68_mem_26_), 
	.A(mem[26]));
   CLKBUF3 FE_PHC67_n726 (.Y(FE_PHN67_n726), 
	.A(n726));
   BUFX2 FE_PHC66_n686 (.Y(FE_PHN66_n686), 
	.A(n686));
   BUFX2 FE_PHC65_FE_OFCN5_n231 (.Y(FE_PHN65_FE_OFCN5_n231), 
	.A(FE_PHN56_FE_OFCN5_n231));
   BUFX2 FE_PHC64_FE_OFCN14_n222 (.Y(FE_PHN64_FE_OFCN14_n222), 
	.A(FE_PHN54_FE_OFCN14_n222));
   BUFX2 FE_PHC63_FE_OFCN12_n224 (.Y(FE_PHN63_FE_OFCN12_n224), 
	.A(FE_OFCN12_n224));
   BUFX2 FE_PHC62_FE_OFCN15_n221 (.Y(FE_PHN62_FE_OFCN15_n221), 
	.A(FE_OFCN15_n221));
   BUFX2 FE_PHC61_FE_OFCN10_n226 (.Y(FE_PHN61_FE_OFCN10_n226), 
	.A(FE_OFCN10_n226));
   BUFX2 FE_PHC60_FE_OFCN7_n229 (.Y(FE_PHN60_FE_OFCN7_n229), 
	.A(FE_OFCN7_n229));
   BUFX2 FE_PHC59_FE_OFCN11_n225 (.Y(FE_PHN59_FE_OFCN11_n225), 
	.A(FE_OFCN11_n225));
   BUFX2 FE_PHC58_FE_OFCN13_n223 (.Y(FE_PHN58_FE_OFCN13_n223), 
	.A(FE_OFCN13_n223));
   BUFX2 FE_PHC57_FE_OFCN8_n228 (.Y(FE_PHN57_FE_OFCN8_n228), 
	.A(FE_OFCN8_n228));
   BUFX2 FE_PHC56_FE_OFCN5_n231 (.Y(FE_PHN56_FE_OFCN5_n231), 
	.A(FE_OFCN5_n231));
   CLKBUF1 FE_PHC55_FE_OFCN16_n219 (.Y(FE_PHN55_FE_OFCN16_n219), 
	.A(FE_OFCN16_n219));
   BUFX2 FE_PHC54_FE_OFCN14_n222 (.Y(FE_PHN54_FE_OFCN14_n222), 
	.A(FE_OFCN14_n222));
   BUFX2 FE_PHC53_FE_OFCN6_n230 (.Y(FE_PHN53_FE_OFCN6_n230), 
	.A(FE_OFCN6_n230));
   CLKBUF1 FE_PHC52_FE_OFCN2_n234 (.Y(FE_PHN52_FE_OFCN2_n234), 
	.A(FE_OFCN2_n234));
   CLKBUF1 FE_PHC51_FE_OFCN4_n232 (.Y(FE_PHN51_FE_OFCN4_n232), 
	.A(FE_OFCN4_n232));
   CLKBUF1 FE_PHC50_FE_OFCN3_n233 (.Y(FE_PHN50_FE_OFCN3_n233), 
	.A(FE_OFCN3_n233));
   CLKBUF1 FE_PHC49_FE_OFCN1_n235 (.Y(FE_PHN49_FE_OFCN1_n235), 
	.A(FE_OFCN1_n235));
   CLKBUF2 FE_PHC48_FE_OFCN9_n227 (.Y(FE_PHN48_FE_OFCN9_n227), 
	.A(FE_OFCN9_n227));
   BUFX2 FE_PSC47_n686 (.Y(FE_PSN47_n686), 
	.A(FE_PHN66_n686));
   BUFX2 FE_PSC46_n34 (.Y(FE_PSN46_n34), 
	.A(n34));
   BUFX2 FE_PSC45_full (.Y(full), 
	.A(FE_PSN45_full));
   BUFX2 FE_PSC44_n36 (.Y(FE_PSN44_n36), 
	.A(n36));
   BUFX2 FE_PSC43_n36 (.Y(FE_PSN43_n36), 
	.A(n36));
   BUFX2 FE_PSC42_FE_OFCN26_n105 (.Y(FE_PSN42_FE_OFCN26_n105), 
	.A(FE_OFCN26_n105));
   BUFX2 FE_PSC41_FE_OFCN28_n123 (.Y(FE_PSN41_FE_OFCN28_n123), 
	.A(FE_OFCN28_n123));
   BUFX4 FE_PSC40_n708 (.Y(FE_PSN40_n708), 
	.A(n708));
   BUFX4 FE_PSC39_FE_OFCN28_n123 (.Y(FE_PSN39_FE_OFCN28_n123), 
	.A(FE_PSN36_FE_OFCN28_n123));
   BUFX4 FE_PSC38_FE_OFCN29_n55 (.Y(FE_PSN38_FE_OFCN29_n55), 
	.A(FE_OFCN29_n55));
   BUFX4 FE_PSC37_n55 (.Y(FE_PSN37_n55), 
	.A(n55));
   BUFX4 FE_PSC36_FE_OFCN28_n123 (.Y(FE_PSN36_FE_OFCN28_n123), 
	.A(FE_OFCN28_n123));
   BUFX4 FE_OFCC29_n55 (.Y(FE_OFCN29_n55), 
	.A(n55));
   BUFX4 FE_OFCC28_n123 (.Y(FE_OFCN28_n123), 
	.A(n123));
   BUFX4 FE_OFCC26_n105 (.Y(FE_OFCN26_n105), 
	.A(n105));
   BUFX4 FE_OFCC20_n199 (.Y(FE_OFCN20_n199), 
	.A(n199));
   BUFX2 FE_OFCC19_n239 (.Y(FE_OFCN19_n239), 
	.A(n239));
   BUFX2 FE_OFCC18_n245 (.Y(FE_OFCN18_n245), 
	.A(n245));
   BUFX4 FE_OFCC17_n241 (.Y(FE_OFCN17_n241), 
	.A(n241));
   BUFX2 FE_OFCC16_n219 (.Y(FE_OFCN16_n219), 
	.A(n219));
   BUFX2 FE_OFCC15_n221 (.Y(FE_OFCN15_n221), 
	.A(n221));
   BUFX2 FE_OFCC14_n222 (.Y(FE_OFCN14_n222), 
	.A(n222));
   BUFX2 FE_OFCC13_n223 (.Y(FE_OFCN13_n223), 
	.A(n223));
   BUFX2 FE_OFCC12_n224 (.Y(FE_OFCN12_n224), 
	.A(n224));
   BUFX2 FE_OFCC11_n225 (.Y(FE_OFCN11_n225), 
	.A(n225));
   BUFX2 FE_OFCC10_n226 (.Y(FE_OFCN10_n226), 
	.A(n226));
   BUFX2 FE_OFCC9_n227 (.Y(FE_OFCN9_n227), 
	.A(n227));
   BUFX2 FE_OFCC8_n228 (.Y(FE_OFCN8_n228), 
	.A(n228));
   BUFX2 FE_OFCC7_n229 (.Y(FE_OFCN7_n229), 
	.A(n229));
   BUFX2 FE_OFCC6_n230 (.Y(FE_OFCN6_n230), 
	.A(n230));
   BUFX2 FE_OFCC5_n231 (.Y(FE_OFCN5_n231), 
	.A(n231));
   BUFX2 FE_OFCC4_n232 (.Y(FE_OFCN4_n232), 
	.A(n232));
   BUFX2 FE_OFCC3_n233 (.Y(FE_OFCN3_n233), 
	.A(n233));
   BUFX2 FE_OFCC2_n234 (.Y(FE_OFCN2_n234), 
	.A(n234));
   BUFX2 FE_OFCC1_n235 (.Y(FE_OFCN1_n235), 
	.A(n235));
   INVX8 clk__L2_I3 (.Y(clk__L2_N3), 
	.A(clk__L1_N0));
   INVX8 clk__L2_I2 (.Y(clk__L2_N2), 
	.A(clk__L1_N0));
   INVX8 clk__L2_I1 (.Y(clk__L2_N1), 
	.A(clk__L1_N0));
   INVX8 clk__L2_I0 (.Y(clk__L2_N0), 
	.A(clk__L1_N0));
   INVX8 clk__L1_I0 (.Y(clk__L1_N0), 
	.A(clk));
   DFFPOSX1 ptr_reg_0_ (.Q(n34), 
	.D(n383), 
	.CLK(clk__L2_N2));
   DFFPOSX1 ptr_reg_1_ (.Q(n35), 
	.D(n381), 
	.CLK(clk__L2_N2));
   DFFPOSX1 empty_reg (.Q(empty), 
	.D(n380), 
	.CLK(clk__L2_N2));
   DFFPOSX1 dout_reg_0_ (.Q(dout[0]), 
	.D(n687), 
	.CLK(clk__L2_N2));
   DFFPOSX1 dout_reg_1_ (.Q(dout[1]), 
	.D(n688), 
	.CLK(clk__L2_N3));
   DFFPOSX1 dout_reg_2_ (.Q(dout[2]), 
	.D(n689), 
	.CLK(clk__L2_N3));
   DFFPOSX1 dout_reg_3_ (.Q(dout[3]), 
	.D(n690), 
	.CLK(clk__L2_N2));
   DFFPOSX1 dout_reg_4_ (.Q(dout[4]), 
	.D(n691), 
	.CLK(clk__L2_N3));
   DFFPOSX1 dout_reg_5_ (.Q(dout[5]), 
	.D(n692), 
	.CLK(clk__L2_N0));
   DFFPOSX1 dout_reg_6_ (.Q(dout[6]), 
	.D(n693), 
	.CLK(clk__L2_N1));
   DFFPOSX1 dout_reg_7_ (.Q(dout[7]), 
	.D(n694), 
	.CLK(clk__L2_N0));
   DFFPOSX1 dout_reg_8_ (.Q(dout[8]), 
	.D(n695), 
	.CLK(clk__L2_N2));
   DFFPOSX1 dout_reg_9_ (.Q(dout[9]), 
	.D(n696), 
	.CLK(clk__L2_N1));
   DFFPOSX1 dout_reg_10_ (.Q(dout[10]), 
	.D(n697), 
	.CLK(clk__L2_N1));
   DFFPOSX1 dout_reg_11_ (.Q(dout[11]), 
	.D(n698), 
	.CLK(clk__L2_N3));
   DFFPOSX1 dout_reg_12_ (.Q(dout[12]), 
	.D(n699), 
	.CLK(clk__L2_N1));
   DFFPOSX1 dout_reg_13_ (.Q(dout[13]), 
	.D(n700), 
	.CLK(clk__L2_N0));
   DFFPOSX1 dout_reg_14_ (.Q(dout[14]), 
	.D(n701), 
	.CLK(clk__L2_N3));
   DFFPOSX1 dout_reg_15_ (.Q(dout[15]), 
	.D(n702), 
	.CLK(clk__L2_N2));
   DFFPOSX1 ptr_reg_2_ (.Q(n36), 
	.D(n382), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_0__15_ (.Q(mem[15]), 
	.D(n364), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_0__14_ (.Q(mem[14]), 
	.D(n365), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_0__13_ (.Q(mem[13]), 
	.D(n366), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_0__12_ (.Q(mem[12]), 
	.D(n367), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_0__11_ (.Q(mem[11]), 
	.D(n368), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_0__10_ (.Q(mem[10]), 
	.D(n369), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_0__9_ (.Q(mem[9]), 
	.D(n370), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_0__8_ (.Q(mem[8]), 
	.D(n371), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_0__7_ (.Q(mem[7]), 
	.D(n372), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_0__6_ (.Q(mem[6]), 
	.D(n373), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_0__5_ (.Q(mem[5]), 
	.D(n374), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_0__4_ (.Q(mem[4]), 
	.D(n375), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_0__3_ (.Q(mem[3]), 
	.D(n376), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_0__2_ (.Q(mem[2]), 
	.D(n377), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_0__1_ (.Q(mem[1]), 
	.D(n378), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_0__0_ (.Q(mem[0]), 
	.D(n379), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_4__15_ (.Q(mem[79]), 
	.D(n300), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__14_ (.Q(mem[78]), 
	.D(n301), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_4__13_ (.Q(mem[77]), 
	.D(n302), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_4__12_ (.Q(mem[76]), 
	.D(n303), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__11_ (.Q(mem[75]), 
	.D(n304), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__10_ (.Q(mem[74]), 
	.D(n305), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__9_ (.Q(mem[73]), 
	.D(n306), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__8_ (.Q(mem[72]), 
	.D(n307), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_4__7_ (.Q(mem[71]), 
	.D(n308), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_4__6_ (.Q(mem[70]), 
	.D(n309), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_4__5_ (.Q(mem[69]), 
	.D(n310), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_4__4_ (.Q(mem[68]), 
	.D(n311), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_4__3_ (.Q(mem[67]), 
	.D(n312), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_4__2_ (.Q(mem[66]), 
	.D(n313), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_4__1_ (.Q(mem[65]), 
	.D(n314), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_4__0_ (.Q(mem[64]), 
	.D(n315), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_1__15_ (.Q(mem[31]), 
	.D(n348), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_1__14_ (.Q(mem[30]), 
	.D(n349), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_1__13_ (.Q(mem[29]), 
	.D(n350), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_1__12_ (.Q(mem[28]), 
	.D(n351), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_1__11_ (.Q(mem[27]), 
	.D(n352), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_1__10_ (.Q(mem[26]), 
	.D(n353), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_1__9_ (.Q(mem[25]), 
	.D(n354), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_1__8_ (.Q(mem[24]), 
	.D(n355), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_1__7_ (.Q(mem[23]), 
	.D(n356), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_1__6_ (.Q(mem[22]), 
	.D(n357), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_1__5_ (.Q(mem[21]), 
	.D(n358), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_1__4_ (.Q(mem[20]), 
	.D(n359), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_1__3_ (.Q(mem[19]), 
	.D(n360), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_1__2_ (.Q(mem[18]), 
	.D(n361), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_1__1_ (.Q(mem[17]), 
	.D(n362), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_1__0_ (.Q(mem[16]), 
	.D(n363), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_2__15_ (.Q(mem[47]), 
	.D(n332), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_2__14_ (.Q(mem[46]), 
	.D(n333), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_2__13_ (.Q(mem[45]), 
	.D(n334), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_2__12_ (.Q(mem[44]), 
	.D(n335), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_2__11_ (.Q(mem[43]), 
	.D(n336), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_2__10_ (.Q(mem[42]), 
	.D(n337), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_2__9_ (.Q(mem[41]), 
	.D(n338), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_2__8_ (.Q(mem[40]), 
	.D(n339), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_2__7_ (.Q(mem[39]), 
	.D(n340), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_2__6_ (.Q(mem[38]), 
	.D(n341), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_2__5_ (.Q(mem[37]), 
	.D(n342), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_2__4_ (.Q(mem[36]), 
	.D(n343), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_2__3_ (.Q(mem[35]), 
	.D(n344), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_2__2_ (.Q(mem[34]), 
	.D(n345), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_2__1_ (.Q(mem[33]), 
	.D(n346), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_2__0_ (.Q(mem[32]), 
	.D(n347), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_6__15_ (.Q(mem[111]), 
	.D(n268), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_6__14_ (.Q(mem[110]), 
	.D(n269), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_6__13_ (.Q(mem[109]), 
	.D(n270), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_6__12_ (.Q(mem[108]), 
	.D(n271), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_6__11_ (.Q(mem[107]), 
	.D(n272), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_6__10_ (.Q(mem[106]), 
	.D(n273), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_6__9_ (.Q(mem[105]), 
	.D(n274), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_6__8_ (.Q(mem[104]), 
	.D(n275), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_6__7_ (.Q(mem[103]), 
	.D(n276), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_6__6_ (.Q(mem[102]), 
	.D(n277), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_6__5_ (.Q(mem[101]), 
	.D(n278), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_6__4_ (.Q(mem[100]), 
	.D(n279), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_6__3_ (.Q(mem[99]), 
	.D(n280), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_6__2_ (.Q(mem[98]), 
	.D(n281), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_6__1_ (.Q(mem[97]), 
	.D(n282), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_6__0_ (.Q(mem[96]), 
	.D(n283), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_7__15_ (.Q(mem[127]), 
	.D(n252), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_7__14_ (.Q(mem[126]), 
	.D(n253), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_7__13_ (.Q(mem[125]), 
	.D(n254), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_7__12_ (.Q(mem[124]), 
	.D(n255), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_7__11_ (.Q(mem[123]), 
	.D(n256), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_7__10_ (.Q(mem[122]), 
	.D(n257), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_7__9_ (.Q(mem[121]), 
	.D(n258), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_7__8_ (.Q(mem[120]), 
	.D(n259), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_7__7_ (.Q(mem[119]), 
	.D(n260), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_7__6_ (.Q(mem[118]), 
	.D(n261), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_7__5_ (.Q(mem[117]), 
	.D(n262), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_7__4_ (.Q(mem[116]), 
	.D(n263), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_7__3_ (.Q(mem[115]), 
	.D(n264), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_7__2_ (.Q(mem[114]), 
	.D(n265), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_7__1_ (.Q(mem[113]), 
	.D(n266), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_7__0_ (.Q(mem[112]), 
	.D(n267), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_3__15_ (.Q(mem[63]), 
	.D(n316), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_3__14_ (.Q(mem[62]), 
	.D(n317), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_3__13_ (.Q(mem[61]), 
	.D(n318), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_3__12_ (.Q(mem[60]), 
	.D(n319), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_3__11_ (.Q(mem[59]), 
	.D(n320), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_3__10_ (.Q(mem[58]), 
	.D(n321), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_3__9_ (.Q(mem[57]), 
	.D(n322), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_3__8_ (.Q(mem[56]), 
	.D(n323), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_3__7_ (.Q(mem[55]), 
	.D(n324), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_3__6_ (.Q(mem[54]), 
	.D(n325), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_3__5_ (.Q(mem[53]), 
	.D(n326), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_3__4_ (.Q(mem[52]), 
	.D(n327), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_3__3_ (.Q(mem[51]), 
	.D(n328), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_3__2_ (.Q(mem[50]), 
	.D(n329), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_3__1_ (.Q(mem[49]), 
	.D(n330), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_3__0_ (.Q(mem[48]), 
	.D(n331), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_5__15_ (.Q(mem[95]), 
	.D(n284), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_5__14_ (.Q(mem[94]), 
	.D(n285), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_5__13_ (.Q(mem[93]), 
	.D(n286), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_5__12_ (.Q(mem[92]), 
	.D(n287), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_5__11_ (.Q(mem[91]), 
	.D(n288), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_5__10_ (.Q(mem[90]), 
	.D(n289), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_5__9_ (.Q(mem[89]), 
	.D(n290), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_5__8_ (.Q(mem[88]), 
	.D(n291), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_5__7_ (.Q(mem[87]), 
	.D(n292), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_5__6_ (.Q(mem[86]), 
	.D(n293), 
	.CLK(clk__L2_N1));
   DFFPOSX1 mem_reg_5__5_ (.Q(mem[85]), 
	.D(n294), 
	.CLK(clk__L2_N0));
   DFFPOSX1 mem_reg_5__4_ (.Q(mem[84]), 
	.D(n295), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_5__3_ (.Q(mem[83]), 
	.D(n296), 
	.CLK(clk__L2_N2));
   DFFPOSX1 mem_reg_5__2_ (.Q(mem[82]), 
	.D(n297), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_5__1_ (.Q(mem[81]), 
	.D(n298), 
	.CLK(clk__L2_N3));
   DFFPOSX1 mem_reg_5__0_ (.Q(mem[80]), 
	.D(n299), 
	.CLK(clk__L2_N0));
   OAI21X1 U55 (.Y(n252), 
	.C(n450), 
	.B(n710), 
	.A(FE_OFCN29_n55));
   OAI21X1 U57 (.Y(n253), 
	.C(n538), 
	.B(n711), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U59 (.Y(n254), 
	.C(n551), 
	.B(n712), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U61 (.Y(n255), 
	.C(n449), 
	.B(n713), 
	.A(FE_PSN37_n55));
   OAI21X1 U63 (.Y(n256), 
	.C(n448), 
	.B(n714), 
	.A(FE_OFCN29_n55));
   OAI21X1 U65 (.Y(n257), 
	.C(n468), 
	.B(n715), 
	.A(FE_PSN37_n55));
   OAI21X1 U67 (.Y(n258), 
	.C(n447), 
	.B(n716), 
	.A(FE_PSN37_n55));
   OAI21X1 U69 (.Y(n259), 
	.C(n446), 
	.B(n717), 
	.A(FE_PSN37_n55));
   OAI21X1 U71 (.Y(n260), 
	.C(n497), 
	.B(n718), 
	.A(FE_OFCN29_n55));
   OAI21X1 U73 (.Y(n261), 
	.C(n506), 
	.B(n719), 
	.A(FE_PSN37_n55));
   OAI21X1 U75 (.Y(n262), 
	.C(n478), 
	.B(n720), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U77 (.Y(n263), 
	.C(n488), 
	.B(n721), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U79 (.Y(n264), 
	.C(n539), 
	.B(n722), 
	.A(FE_OFCN29_n55));
   OAI21X1 U81 (.Y(n265), 
	.C(n552), 
	.B(n723), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U83 (.Y(n266), 
	.C(n515), 
	.B(n724), 
	.A(FE_PSN38_FE_OFCN29_n55));
   OAI21X1 U85 (.Y(n267), 
	.C(n526), 
	.B(n725), 
	.A(FE_OFCN29_n55));
   NAND3X1 U87 (.Y(n55), 
	.C(n707), 
	.B(FE_PSN44_n36), 
	.A(n179));
   OAI21X1 U88 (.Y(n268), 
	.C(n536), 
	.B(n684), 
	.A(n710));
   OAI21X1 U90 (.Y(n269), 
	.C(n549), 
	.B(n684), 
	.A(n711));
   OAI21X1 U92 (.Y(n270), 
	.C(n445), 
	.B(n684), 
	.A(n712));
   OAI21X1 U94 (.Y(n271), 
	.C(n444), 
	.B(n684), 
	.A(n713));
   OAI21X1 U96 (.Y(n272), 
	.C(n467), 
	.B(n684), 
	.A(n714));
   OAI21X1 U98 (.Y(n273), 
	.C(n443), 
	.B(n684), 
	.A(n715));
   OAI21X1 U100 (.Y(n274), 
	.C(n442), 
	.B(n684), 
	.A(n716));
   OAI21X1 U102 (.Y(n275), 
	.C(n441), 
	.B(n684), 
	.A(n717));
   OAI21X1 U104 (.Y(n276), 
	.C(n505), 
	.B(n684), 
	.A(n718));
   OAI21X1 U106 (.Y(n277), 
	.C(n496), 
	.B(n684), 
	.A(n719));
   OAI21X1 U108 (.Y(n278), 
	.C(n487), 
	.B(n684), 
	.A(n720));
   OAI21X1 U110 (.Y(n279), 
	.C(n477), 
	.B(n684), 
	.A(n721));
   OAI21X1 U112 (.Y(n280), 
	.C(n550), 
	.B(n684), 
	.A(n722));
   OAI21X1 U114 (.Y(n281), 
	.C(n537), 
	.B(n684), 
	.A(n723));
   OAI21X1 U116 (.Y(n282), 
	.C(n525), 
	.B(n684), 
	.A(n724));
   OAI21X1 U118 (.Y(n283), 
	.C(n514), 
	.B(n684), 
	.A(n725));
   OAI21X1 U121 (.Y(n284), 
	.C(n518), 
	.B(FE_OFCN26_n105), 
	.A(n710));
   OAI21X1 U123 (.Y(n285), 
	.C(n529), 
	.B(FE_OFCN26_n105), 
	.A(n711));
   OAI21X1 U125 (.Y(n286), 
	.C(n440), 
	.B(FE_OFCN26_n105), 
	.A(n712));
   OAI21X1 U127 (.Y(n287), 
	.C(n439), 
	.B(FE_OFCN26_n105), 
	.A(n713));
   OAI21X1 U129 (.Y(n288), 
	.C(n438), 
	.B(FE_OFCN26_n105), 
	.A(n714));
   OAI21X1 U131 (.Y(n289), 
	.C(n437), 
	.B(FE_OFCN26_n105), 
	.A(n715));
   OAI21X1 U133 (.Y(n290), 
	.C(n436), 
	.B(FE_OFCN26_n105), 
	.A(n716));
   OAI21X1 U135 (.Y(n291), 
	.C(n470), 
	.B(FE_OFCN26_n105), 
	.A(n717));
   OAI21X1 U137 (.Y(n292), 
	.C(n480), 
	.B(FE_PSN42_FE_OFCN26_n105), 
	.A(n718));
   OAI21X1 U139 (.Y(n293), 
	.C(n490), 
	.B(FE_OFCN26_n105), 
	.A(n719));
   OAI21X1 U141 (.Y(n294), 
	.C(n499), 
	.B(FE_OFCN26_n105), 
	.A(n720));
   OAI21X1 U143 (.Y(n295), 
	.C(n508), 
	.B(FE_OFCN26_n105), 
	.A(n721));
   OAI21X1 U145 (.Y(n296), 
	.C(n519), 
	.B(FE_OFCN26_n105), 
	.A(n722));
   OAI21X1 U147 (.Y(n297), 
	.C(n530), 
	.B(FE_OFCN26_n105), 
	.A(n723));
   OAI21X1 U149 (.Y(n298), 
	.C(n541), 
	.B(FE_OFCN26_n105), 
	.A(n724));
   OAI21X1 U151 (.Y(n299), 
	.C(n554), 
	.B(FE_PSN42_FE_OFCN26_n105), 
	.A(n725));
   NAND3X1 U153 (.Y(n105), 
	.C(FE_PSN44_n36), 
	.B(n685), 
	.A(n705));
   OAI21X1 U154 (.Y(n300), 
	.C(n435), 
	.B(n710), 
	.A(FE_OFCN28_n123));
   OAI21X1 U156 (.Y(n301), 
	.C(n464), 
	.B(n711), 
	.A(FE_PSN39_FE_OFCN28_n123));
   OAI21X1 U158 (.Y(n302), 
	.C(n510), 
	.B(n712), 
	.A(FE_PSN39_FE_OFCN28_n123));
   OAI21X1 U160 (.Y(n303), 
	.C(n521), 
	.B(n713), 
	.A(FE_OFCN28_n123));
   OAI21X1 U162 (.Y(n304), 
	.C(n532), 
	.B(n714), 
	.A(FE_OFCN28_n123));
   OAI21X1 U164 (.Y(n305), 
	.C(n545), 
	.B(n715), 
	.A(FE_OFCN28_n123));
   OAI21X1 U166 (.Y(n306), 
	.C(n434), 
	.B(n716), 
	.A(FE_OFCN28_n123));
   OAI21X1 U168 (.Y(n307), 
	.C(n433), 
	.B(n717), 
	.A(n123));
   OAI21X1 U170 (.Y(n308), 
	.C(n533), 
	.B(n718), 
	.A(FE_PSN39_FE_OFCN28_n123));
   OAI21X1 U172 (.Y(n309), 
	.C(n546), 
	.B(n719), 
	.A(n123));
   OAI21X1 U174 (.Y(n310), 
	.C(n511), 
	.B(n720), 
	.A(FE_PSN39_FE_OFCN28_n123));
   OAI21X1 U176 (.Y(n311), 
	.C(n522), 
	.B(n721), 
	.A(FE_PSN39_FE_OFCN28_n123));
   OAI21X1 U178 (.Y(n312), 
	.C(n493), 
	.B(n722), 
	.A(n123));
   OAI21X1 U180 (.Y(n313), 
	.C(n502), 
	.B(n723), 
	.A(FE_PSN41_FE_OFCN28_n123));
   OAI21X1 U182 (.Y(n314), 
	.C(n472), 
	.B(n724), 
	.A(FE_OFCN28_n123));
   OAI21X1 U184 (.Y(n315), 
	.C(n482), 
	.B(n725), 
	.A(FE_PSN39_FE_OFCN28_n123));
   NAND3X1 U186 (.Y(n141), 
	.C(n160), 
	.B(FE_PSN46_n34), 
	.A(n707));
   NAND3X1 U187 (.Y(n140), 
	.C(n248), 
	.B(FE_PSN44_n36), 
	.A(n706));
   OAI21X1 U188 (.Y(n316), 
	.C(n527), 
	.B(n683), 
	.A(n710));
   OAI21X1 U190 (.Y(n317), 
	.C(n516), 
	.B(n683), 
	.A(n711));
   OAI21X1 U192 (.Y(n318), 
	.C(n432), 
	.B(n683), 
	.A(n712));
   OAI21X1 U194 (.Y(n319), 
	.C(n431), 
	.B(n683), 
	.A(n713));
   OAI21X1 U196 (.Y(n320), 
	.C(n430), 
	.B(n683), 
	.A(n714));
   OAI21X1 U198 (.Y(n321), 
	.C(n429), 
	.B(n683), 
	.A(n715));
   OAI21X1 U200 (.Y(n322), 
	.C(n469), 
	.B(n683), 
	.A(n716));
   OAI21X1 U202 (.Y(n323), 
	.C(n428), 
	.B(n683), 
	.A(n717));
   OAI21X1 U204 (.Y(n324), 
	.C(n489), 
	.B(n683), 
	.A(n718));
   OAI21X1 U206 (.Y(n325), 
	.C(n479), 
	.B(n683), 
	.A(n719));
   OAI21X1 U208 (.Y(n326), 
	.C(n507), 
	.B(n683), 
	.A(n720));
   OAI21X1 U210 (.Y(n327), 
	.C(n498), 
	.B(n683), 
	.A(n721));
   OAI21X1 U212 (.Y(n328), 
	.C(n528), 
	.B(n683), 
	.A(n722));
   OAI21X1 U214 (.Y(n329), 
	.C(n517), 
	.B(n683), 
	.A(n723));
   OAI21X1 U216 (.Y(n330), 
	.C(n553), 
	.B(n683), 
	.A(n724));
   OAI21X1 U218 (.Y(n331), 
	.C(n540), 
	.B(n683), 
	.A(n725));
   AOI22X1 U221 (.Y(n159), 
	.D(FE_PSN46_n34), 
	.C(n706), 
	.B(n686), 
	.A(n707));
   OAI21X1 U222 (.Y(n332), 
	.C(n475), 
	.B(n682), 
	.A(n710));
   OAI21X1 U224 (.Y(n333), 
	.C(n485), 
	.B(n682), 
	.A(n711));
   OAI21X1 U226 (.Y(n334), 
	.C(n427), 
	.B(n682), 
	.A(n712));
   OAI21X1 U228 (.Y(n335), 
	.C(n466), 
	.B(n682), 
	.A(n713));
   OAI21X1 U230 (.Y(n336), 
	.C(n426), 
	.B(n682), 
	.A(n714));
   OAI21X1 U232 (.Y(n337), 
	.C(n425), 
	.B(n682), 
	.A(n715));
   OAI21X1 U234 (.Y(n338), 
	.C(n424), 
	.B(n682), 
	.A(n716));
   OAI21X1 U236 (.Y(n339), 
	.C(n423), 
	.B(n682), 
	.A(n717));
   OAI21X1 U238 (.Y(n340), 
	.C(n513), 
	.B(n682), 
	.A(n718));
   OAI21X1 U240 (.Y(n341), 
	.C(n524), 
	.B(n682), 
	.A(n719));
   OAI21X1 U242 (.Y(n342), 
	.C(n535), 
	.B(n682), 
	.A(n720));
   OAI21X1 U244 (.Y(n343), 
	.C(n548), 
	.B(n682), 
	.A(n721));
   OAI21X1 U246 (.Y(n344), 
	.C(n476), 
	.B(n682), 
	.A(n722));
   OAI21X1 U248 (.Y(n345), 
	.C(n486), 
	.B(n682), 
	.A(n723));
   OAI21X1 U250 (.Y(n346), 
	.C(n495), 
	.B(n682), 
	.A(n724));
   OAI21X1 U252 (.Y(n347), 
	.C(n504), 
	.B(n682), 
	.A(n725));
   AOI22X1 U255 (.Y(n178), 
	.D(n179), 
	.C(n706), 
	.B(n707), 
	.A(n180));
   OAI21X1 U256 (.Y(n348), 
	.C(n465), 
	.B(n710), 
	.A(n181));
   OAI21X1 U258 (.Y(n349), 
	.C(n473), 
	.B(n711), 
	.A(n181));
   OAI21X1 U260 (.Y(n350), 
	.C(n483), 
	.B(n712), 
	.A(n181));
   OAI21X1 U262 (.Y(n351), 
	.C(n422), 
	.B(n713), 
	.A(n181));
   OAI21X1 U264 (.Y(n352), 
	.C(n421), 
	.B(n714), 
	.A(n181));
   OAI21X1 U266 (.Y(n353), 
	.C(n420), 
	.B(n715), 
	.A(n181));
   OAI21X1 U268 (.Y(n354), 
	.C(n419), 
	.B(n716), 
	.A(n181));
   OAI21X1 U270 (.Y(n355), 
	.C(n418), 
	.B(n717), 
	.A(n181));
   OAI21X1 U272 (.Y(n356), 
	.C(n523), 
	.B(n718), 
	.A(n181));
   OAI21X1 U274 (.Y(n357), 
	.C(n512), 
	.B(n719), 
	.A(n181));
   OAI21X1 U276 (.Y(n358), 
	.C(n547), 
	.B(n720), 
	.A(n181));
   OAI21X1 U278 (.Y(n359), 
	.C(n534), 
	.B(n721), 
	.A(n181));
   OAI21X1 U280 (.Y(n360), 
	.C(n484), 
	.B(n722), 
	.A(n181));
   OAI21X1 U282 (.Y(n361), 
	.C(n474), 
	.B(n723), 
	.A(n181));
   OAI21X1 U284 (.Y(n362), 
	.C(n503), 
	.B(n724), 
	.A(n181));
   OAI21X1 U286 (.Y(n363), 
	.C(n494), 
	.B(n725), 
	.A(n181));
   AOI21X1 U288 (.Y(n181), 
	.C(n198), 
	.B(n237), 
	.A(n707));
   NOR3X1 U289 (.Y(n198), 
	.C(FE_OFCN20_n199), 
	.B(FE_PSN44_n36), 
	.A(n557));
   NAND3X1 U290 (.Y(n200), 
	.C(n201), 
	.B(n709), 
	.A(n726));
   OAI21X1 U291 (.Y(n364), 
	.C(n491), 
	.B(n681), 
	.A(n710));
   OAI21X1 U293 (.Y(n365), 
	.C(n500), 
	.B(n681), 
	.A(n711));
   OAI21X1 U295 (.Y(n366), 
	.C(n463), 
	.B(n681), 
	.A(n712));
   OAI21X1 U297 (.Y(n367), 
	.C(n417), 
	.B(n681), 
	.A(n713));
   OAI21X1 U299 (.Y(n368), 
	.C(n416), 
	.B(n681), 
	.A(n714));
   OAI21X1 U301 (.Y(n369), 
	.C(n415), 
	.B(n681), 
	.A(n715));
   OAI21X1 U303 (.Y(n370), 
	.C(n414), 
	.B(n681), 
	.A(n716));
   OAI21X1 U305 (.Y(n371), 
	.C(n413), 
	.B(n681), 
	.A(n717));
   OAI21X1 U307 (.Y(n372), 
	.C(n544), 
	.B(n681), 
	.A(n718));
   OAI21X1 U309 (.Y(n373), 
	.C(n531), 
	.B(n681), 
	.A(n719));
   OAI21X1 U311 (.Y(n374), 
	.C(n520), 
	.B(n681), 
	.A(n720));
   OAI21X1 U313 (.Y(n375), 
	.C(n509), 
	.B(n681), 
	.A(n721));
   OAI21X1 U315 (.Y(n376), 
	.C(n501), 
	.B(n681), 
	.A(n722));
   OAI21X1 U317 (.Y(n377), 
	.C(n492), 
	.B(n681), 
	.A(n723));
   OAI21X1 U319 (.Y(n378), 
	.C(n481), 
	.B(n681), 
	.A(n724));
   OAI21X1 U321 (.Y(n379), 
	.C(n471), 
	.B(n681), 
	.A(n725));
   NAND3X1 U324 (.Y(n199), 
	.C(empty), 
	.B(n709), 
	.A(n201));
   AOI22X1 U325 (.Y(n219), 
	.D(n220), 
	.C(n64), 
	.B(n555), 
	.A(dout[15]));
   AOI22X1 U326 (.Y(n221), 
	.D(n220), 
	.C(n65), 
	.B(n555), 
	.A(dout[14]));
   AOI22X1 U327 (.Y(n222), 
	.D(n220), 
	.C(n66), 
	.B(n555), 
	.A(dout[13]));
   AOI22X1 U328 (.Y(n223), 
	.D(n220), 
	.C(n67), 
	.B(n555), 
	.A(dout[12]));
   AOI22X1 U329 (.Y(n224), 
	.D(n220), 
	.C(n68), 
	.B(n555), 
	.A(dout[11]));
   AOI22X1 U330 (.Y(n225), 
	.D(n220), 
	.C(n69), 
	.B(n555), 
	.A(dout[10]));
   AOI22X1 U331 (.Y(n226), 
	.D(n220), 
	.C(n70), 
	.B(n555), 
	.A(dout[9]));
   AOI22X1 U332 (.Y(n227), 
	.D(n220), 
	.C(n71), 
	.B(n555), 
	.A(dout[8]));
   AOI22X1 U333 (.Y(n228), 
	.D(n220), 
	.C(n72), 
	.B(n555), 
	.A(dout[7]));
   AOI22X1 U334 (.Y(n229), 
	.D(n220), 
	.C(n73), 
	.B(n555), 
	.A(dout[6]));
   AOI22X1 U335 (.Y(n230), 
	.D(n220), 
	.C(n74), 
	.B(n555), 
	.A(dout[5]));
   AOI22X1 U336 (.Y(n231), 
	.D(n220), 
	.C(n75), 
	.B(n555), 
	.A(dout[4]));
   AOI22X1 U337 (.Y(n232), 
	.D(n220), 
	.C(n76), 
	.B(n555), 
	.A(dout[3]));
   AOI22X1 U338 (.Y(n233), 
	.D(n220), 
	.C(n77), 
	.B(n555), 
	.A(dout[2]));
   AOI22X1 U339 (.Y(n234), 
	.D(n220), 
	.C(n78), 
	.B(n555), 
	.A(dout[1]));
   AOI22X1 U340 (.Y(n235), 
	.D(n220), 
	.C(n79), 
	.B(n555), 
	.A(dout[0]));
   OAI21X1 U341 (.Y(n380), 
	.C(n236), 
	.B(FE_PHN67_n726), 
	.A(n201));
   AOI21X1 U342 (.Y(n236), 
	.C(reset), 
	.B(n237), 
	.A(n703));
   NAND3X1 U343 (.Y(n381), 
	.C(n455), 
	.B(FE_OFCN19_n239), 
	.A(n238));
   NAND3X1 U345 (.Y(n239), 
	.C(n242), 
	.B(FE_OFCN17_n241), 
	.A(n220));
   NAND3X1 U346 (.Y(n238), 
	.C(n462), 
	.B(n458), 
	.A(n461));
   OAI21X1 U350 (.Y(n382), 
	.C(n246), 
	.B(n727), 
	.A(FE_OFCN18_n245));
   NAND3X1 U351 (.Y(n246), 
	.C(n462), 
	.B(n461), 
	.A(FE_PHN74_n247));
   OAI21X1 U352 (.Y(n247), 
	.C(n727), 
	.B(n556), 
	.A(FE_PSN47_n686));
   AOI21X1 U354 (.Y(n245), 
	.C(n459), 
	.B(n542), 
	.A(n220));
   OAI21X1 U356 (.Y(n383), 
	.C(n412), 
	.B(FE_OFCN17_n241), 
	.A(FE_PSN47_n686));
   NAND3X1 U359 (.Y(n241), 
	.C(n454), 
	.B(n709), 
	.A(n461));
   NOR3X1 U361 (.Y(n201), 
	.C(n708), 
	.B(pop), 
	.A(FE_PSN45_full));
   NAND3X1 U365 (.Y(n251), 
	.C(pop), 
	.B(FE_PSN40_n708), 
	.A(n726));
   NOR3X1 U366 (.Y(FE_PSN45_full), 
	.C(n727), 
	.B(n686), 
	.A(n685));
   AND2X1 U367 (.Y(n243), 
	.B(n457), 
	.A(n703));
   AND2X2 U368 (.Y(n123), 
	.B(n141), 
	.A(n140));
   AND2X2 U369 (.Y(n242), 
	.B(n557), 
	.A(n456));
   AND2X2 U398 (.Y(n249), 
	.B(FE_PSN47_n686), 
	.A(n462));
   INVX1 U399 (.Y(n412), 
	.A(n249));
   AND2X1 U400 (.Y(n210), 
	.B(n681), 
	.A(mem[8]));
   INVX1 U401 (.Y(n413), 
	.A(n210));
   AND2X1 U402 (.Y(n209), 
	.B(n681), 
	.A(mem[9]));
   INVX1 U403 (.Y(n414), 
	.A(n209));
   AND2X1 U404 (.Y(n208), 
	.B(n681), 
	.A(mem[10]));
   INVX1 U405 (.Y(n415), 
	.A(n208));
   AND2X1 U406 (.Y(n207), 
	.B(n681), 
	.A(mem[11]));
   INVX1 U407 (.Y(n416), 
	.A(n207));
   AND2X1 U408 (.Y(n206), 
	.B(n681), 
	.A(mem[12]));
   INVX1 U409 (.Y(n417), 
	.A(n206));
   AND2X1 U410 (.Y(n189), 
	.B(n181), 
	.A(mem[24]));
   INVX1 U411 (.Y(n418), 
	.A(n189));
   AND2X1 U412 (.Y(n188), 
	.B(n181), 
	.A(mem[25]));
   INVX1 U413 (.Y(n419), 
	.A(n188));
   AND2X1 U414 (.Y(n187), 
	.B(n181), 
	.A(FE_PHN68_mem_26_));
   INVX1 U415 (.Y(n420), 
	.A(n187));
   AND2X2 U416 (.Y(n186), 
	.B(n181), 
	.A(FE_PHN78_mem_27_));
   INVX2 U417 (.Y(n421), 
	.A(n186));
   AND2X2 U418 (.Y(n185), 
	.B(n181), 
	.A(FE_PHN73_mem_28_));
   INVX2 U419 (.Y(n422), 
	.A(n185));
   AND2X1 U420 (.Y(n169), 
	.B(n682), 
	.A(mem[40]));
   INVX1 U421 (.Y(n423), 
	.A(n169));
   AND2X1 U422 (.Y(n168), 
	.B(n682), 
	.A(mem[41]));
   INVX1 U423 (.Y(n424), 
	.A(n168));
   AND2X1 U424 (.Y(n167), 
	.B(n682), 
	.A(mem[42]));
   INVX1 U425 (.Y(n425), 
	.A(n167));
   AND2X1 U426 (.Y(n166), 
	.B(n682), 
	.A(mem[43]));
   INVX1 U427 (.Y(n426), 
	.A(n166));
   AND2X1 U428 (.Y(n164), 
	.B(n682), 
	.A(mem[45]));
   INVX1 U429 (.Y(n427), 
	.A(n164));
   AND2X1 U430 (.Y(n150), 
	.B(n683), 
	.A(mem[56]));
   INVX1 U431 (.Y(n428), 
	.A(n150));
   AND2X1 U432 (.Y(n148), 
	.B(n683), 
	.A(mem[58]));
   INVX1 U433 (.Y(n429), 
	.A(n148));
   AND2X1 U434 (.Y(n147), 
	.B(n683), 
	.A(mem[59]));
   INVX1 U435 (.Y(n430), 
	.A(n147));
   AND2X1 U436 (.Y(n146), 
	.B(n683), 
	.A(mem[60]));
   INVX1 U437 (.Y(n431), 
	.A(n146));
   AND2X1 U438 (.Y(n145), 
	.B(n683), 
	.A(mem[61]));
   INVX1 U439 (.Y(n432), 
	.A(n145));
   AND2X2 U440 (.Y(n131), 
	.B(n123), 
	.A(mem[72]));
   INVX1 U441 (.Y(n433), 
	.A(n131));
   AND2X1 U442 (.Y(n130), 
	.B(FE_OFCN28_n123), 
	.A(mem[73]));
   INVX1 U443 (.Y(n434), 
	.A(n130));
   AND2X1 U444 (.Y(n124), 
	.B(FE_OFCN28_n123), 
	.A(mem[79]));
   INVX1 U445 (.Y(n435), 
	.A(n124));
   AND2X1 U446 (.Y(n112), 
	.B(FE_OFCN26_n105), 
	.A(mem[89]));
   INVX1 U447 (.Y(n436), 
	.A(n112));
   AND2X1 U448 (.Y(n111), 
	.B(FE_OFCN26_n105), 
	.A(mem[90]));
   INVX1 U449 (.Y(n437), 
	.A(n111));
   AND2X1 U450 (.Y(n110), 
	.B(FE_OFCN26_n105), 
	.A(mem[91]));
   INVX1 U451 (.Y(n438), 
	.A(n110));
   AND2X1 U452 (.Y(n109), 
	.B(FE_OFCN26_n105), 
	.A(mem[92]));
   INVX1 U453 (.Y(n439), 
	.A(n109));
   AND2X1 U454 (.Y(n108), 
	.B(FE_OFCN26_n105), 
	.A(mem[93]));
   INVX1 U455 (.Y(n440), 
	.A(n108));
   AND2X1 U456 (.Y(n96), 
	.B(n684), 
	.A(mem[104]));
   INVX1 U457 (.Y(n441), 
	.A(n96));
   AND2X1 U458 (.Y(n95), 
	.B(n684), 
	.A(mem[105]));
   INVX1 U459 (.Y(n442), 
	.A(n95));
   AND2X1 U460 (.Y(n94), 
	.B(n684), 
	.A(mem[106]));
   INVX1 U461 (.Y(n443), 
	.A(n94));
   AND2X1 U462 (.Y(n92), 
	.B(n684), 
	.A(mem[108]));
   INVX1 U463 (.Y(n444), 
	.A(n92));
   AND2X1 U464 (.Y(n91), 
	.B(n684), 
	.A(mem[109]));
   INVX1 U465 (.Y(n445), 
	.A(n91));
   AND2X2 U466 (.Y(n63), 
	.B(FE_PSN37_n55), 
	.A(mem[120]));
   INVX1 U467 (.Y(n446), 
	.A(n63));
   AND2X2 U468 (.Y(n62), 
	.B(FE_PSN37_n55), 
	.A(mem[121]));
   INVX1 U469 (.Y(n447), 
	.A(n62));
   AND2X1 U470 (.Y(n60), 
	.B(FE_OFCN29_n55), 
	.A(mem[123]));
   INVX1 U471 (.Y(n448), 
	.A(n60));
   AND2X1 U472 (.Y(n59), 
	.B(FE_PSN37_n55), 
	.A(mem[124]));
   INVX1 U473 (.Y(n449), 
	.A(n59));
   AND2X2 U474 (.Y(n56), 
	.B(FE_OFCN29_n55), 
	.A(mem[127]));
   INVX1 U475 (.Y(n450), 
	.A(n56));
   AND2X1 U479 (.Y(n250), 
	.B(n726), 
	.A(n201));
   INVX2 U480 (.Y(n454), 
	.A(n250));
   AND2X1 U481 (.Y(n240), 
	.B(n678), 
	.A(n459));
   INVX1 U482 (.Y(n455), 
	.A(n240));
   AND2X1 U483 (.Y(n179), 
	.B(n686), 
	.A(n678));
   INVX1 U484 (.Y(n456), 
	.A(n179));
   AND2X1 U485 (.Y(n237), 
	.B(n727), 
	.A(n248));
   INVX1 U486 (.Y(n457), 
	.A(n237));
   INVX2 U487 (.Y(n458), 
	.A(n242));
   INVX2 U488 (.Y(n459), 
	.A(FE_OFCN17_n241));
   INVX2 U490 (.Y(n461), 
	.A(n243));
   OR2X2 U491 (.Y(n244), 
	.B(reset), 
	.A(n459));
   INVX4 U492 (.Y(n462), 
	.A(n244));
   AND2X1 U493 (.Y(n205), 
	.B(n681), 
	.A(mem[13]));
   INVX1 U494 (.Y(n463), 
	.A(n205));
   AND2X1 U495 (.Y(n125), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(mem[78]));
   INVX1 U496 (.Y(n464), 
	.A(n125));
   AND2X1 U497 (.Y(n182), 
	.B(n181), 
	.A(FE_PHN77_mem_31_));
   INVX1 U498 (.Y(n465), 
	.A(n182));
   AND2X1 U499 (.Y(n165), 
	.B(n682), 
	.A(mem[44]));
   INVX1 U500 (.Y(n466), 
	.A(n165));
   AND2X1 U501 (.Y(n93), 
	.B(n684), 
	.A(mem[107]));
   INVX1 U502 (.Y(n467), 
	.A(n93));
   AND2X2 U503 (.Y(n61), 
	.B(FE_PSN37_n55), 
	.A(mem[122]));
   INVX1 U504 (.Y(n468), 
	.A(n61));
   AND2X1 U505 (.Y(n149), 
	.B(n683), 
	.A(mem[57]));
   INVX1 U506 (.Y(n469), 
	.A(n149));
   AND2X1 U507 (.Y(n114), 
	.B(n105), 
	.A(mem[88]));
   INVX1 U508 (.Y(n470), 
	.A(n114));
   AND2X1 U509 (.Y(n218), 
	.B(n681), 
	.A(mem[0]));
   INVX1 U510 (.Y(n471), 
	.A(n218));
   AND2X2 U511 (.Y(n138), 
	.B(FE_PSN36_FE_OFCN28_n123), 
	.A(mem[65]));
   INVX1 U512 (.Y(n472), 
	.A(n138));
   AND2X1 U513 (.Y(n183), 
	.B(n181), 
	.A(FE_PHN71_mem_30_));
   INVX1 U514 (.Y(n473), 
	.A(n183));
   AND2X1 U515 (.Y(n195), 
	.B(n181), 
	.A(mem[18]));
   INVX1 U516 (.Y(n474), 
	.A(n195));
   AND2X1 U517 (.Y(n162), 
	.B(n682), 
	.A(FE_PHN81_mem_47_));
   INVX1 U518 (.Y(n475), 
	.A(n162));
   AND2X1 U519 (.Y(n174), 
	.B(n682), 
	.A(mem[35]));
   INVX1 U520 (.Y(n476), 
	.A(n174));
   AND2X1 U521 (.Y(n100), 
	.B(n684), 
	.A(mem[100]));
   INVX1 U522 (.Y(n477), 
	.A(n100));
   AND2X2 U523 (.Y(n82), 
	.B(FE_PSN38_FE_OFCN29_n55), 
	.A(mem[117]));
   INVX1 U524 (.Y(n478), 
	.A(n82));
   AND2X1 U525 (.Y(n152), 
	.B(n683), 
	.A(mem[54]));
   INVX1 U526 (.Y(n479), 
	.A(n152));
   AND2X1 U527 (.Y(n115), 
	.B(FE_OFCN26_n105), 
	.A(mem[87]));
   INVX1 U528 (.Y(n480), 
	.A(n115));
   AND2X1 U529 (.Y(n217), 
	.B(n681), 
	.A(mem[1]));
   INVX1 U530 (.Y(n481), 
	.A(n217));
   AND2X2 U531 (.Y(n139), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(mem[64]));
   INVX1 U532 (.Y(n482), 
	.A(n139));
   AND2X1 U533 (.Y(n184), 
	.B(n181), 
	.A(FE_PHN70_mem_29_));
   INVX1 U534 (.Y(n483), 
	.A(n184));
   AND2X1 U535 (.Y(n194), 
	.B(n181), 
	.A(FE_PHN76_mem_19_));
   INVX2 U536 (.Y(n484), 
	.A(n194));
   AND2X1 U537 (.Y(n163), 
	.B(n682), 
	.A(mem[46]));
   INVX1 U538 (.Y(n485), 
	.A(n163));
   AND2X1 U539 (.Y(n175), 
	.B(n682), 
	.A(mem[34]));
   INVX1 U540 (.Y(n486), 
	.A(n175));
   AND2X1 U541 (.Y(n99), 
	.B(n684), 
	.A(mem[101]));
   INVX1 U542 (.Y(n487), 
	.A(n99));
   AND2X1 U543 (.Y(n83), 
	.B(FE_PSN38_FE_OFCN29_n55), 
	.A(mem[116]));
   INVX1 U544 (.Y(n488), 
	.A(n83));
   AND2X1 U545 (.Y(n151), 
	.B(n683), 
	.A(mem[55]));
   INVX1 U546 (.Y(n489), 
	.A(n151));
   AND2X1 U547 (.Y(n116), 
	.B(FE_OFCN26_n105), 
	.A(mem[86]));
   INVX1 U548 (.Y(n490), 
	.A(n116));
   AND2X1 U549 (.Y(n203), 
	.B(n681), 
	.A(mem[15]));
   INVX1 U550 (.Y(n491), 
	.A(n203));
   AND2X1 U551 (.Y(n216), 
	.B(n681), 
	.A(mem[2]));
   INVX1 U552 (.Y(n492), 
	.A(n216));
   AND2X2 U553 (.Y(n136), 
	.B(n123), 
	.A(mem[67]));
   INVX1 U554 (.Y(n493), 
	.A(n136));
   AND2X1 U555 (.Y(n197), 
	.B(n181), 
	.A(FE_PHN82_mem_16_));
   INVX1 U556 (.Y(n494), 
	.A(n197));
   AND2X1 U557 (.Y(n176), 
	.B(n682), 
	.A(mem[33]));
   INVX1 U558 (.Y(n495), 
	.A(n176));
   AND2X1 U559 (.Y(n98), 
	.B(n684), 
	.A(mem[102]));
   INVX1 U560 (.Y(n496), 
	.A(n98));
   AND2X1 U561 (.Y(n80), 
	.B(FE_OFCN29_n55), 
	.A(FE_PHN79_mem_119_));
   INVX1 U562 (.Y(n497), 
	.A(n80));
   AND2X1 U563 (.Y(n154), 
	.B(n683), 
	.A(mem[52]));
   INVX1 U564 (.Y(n498), 
	.A(n154));
   AND2X1 U565 (.Y(n117), 
	.B(FE_OFCN26_n105), 
	.A(mem[85]));
   INVX1 U566 (.Y(n499), 
	.A(n117));
   AND2X1 U567 (.Y(n204), 
	.B(n681), 
	.A(mem[14]));
   INVX1 U568 (.Y(n500), 
	.A(n204));
   AND2X1 U569 (.Y(n215), 
	.B(n681), 
	.A(mem[3]));
   INVX1 U570 (.Y(n501), 
	.A(n215));
   AND2X2 U571 (.Y(n137), 
	.B(FE_OFCN28_n123), 
	.A(mem[66]));
   INVX1 U572 (.Y(n502), 
	.A(n137));
   AND2X1 U573 (.Y(n196), 
	.B(n181), 
	.A(mem[17]));
   INVX1 U574 (.Y(n503), 
	.A(n196));
   AND2X1 U575 (.Y(n177), 
	.B(n682), 
	.A(mem[32]));
   INVX1 U576 (.Y(n504), 
	.A(n177));
   AND2X1 U577 (.Y(n97), 
	.B(n684), 
	.A(mem[103]));
   INVX1 U578 (.Y(n505), 
	.A(n97));
   AND2X1 U579 (.Y(n81), 
	.B(FE_PSN37_n55), 
	.A(mem[118]));
   INVX1 U580 (.Y(n506), 
	.A(n81));
   AND2X1 U581 (.Y(n153), 
	.B(n683), 
	.A(mem[53]));
   INVX1 U582 (.Y(n507), 
	.A(n153));
   AND2X1 U583 (.Y(n118), 
	.B(FE_OFCN26_n105), 
	.A(mem[84]));
   INVX1 U584 (.Y(n508), 
	.A(n118));
   AND2X1 U585 (.Y(n214), 
	.B(n681), 
	.A(mem[4]));
   INVX1 U586 (.Y(n509), 
	.A(n214));
   AND2X2 U587 (.Y(n126), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(mem[77]));
   INVX1 U588 (.Y(n510), 
	.A(n126));
   AND2X1 U589 (.Y(n134), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(mem[69]));
   INVX1 U590 (.Y(n511), 
	.A(n134));
   AND2X1 U591 (.Y(n191), 
	.B(n181), 
	.A(mem[22]));
   INVX1 U592 (.Y(n512), 
	.A(n191));
   AND2X1 U593 (.Y(n170), 
	.B(n682), 
	.A(mem[39]));
   INVX1 U594 (.Y(n513), 
	.A(n170));
   AND2X1 U595 (.Y(n104), 
	.B(n684), 
	.A(mem[96]));
   INVX1 U596 (.Y(n514), 
	.A(n104));
   AND2X2 U597 (.Y(n86), 
	.B(FE_PSN38_FE_OFCN29_n55), 
	.A(mem[113]));
   INVX1 U598 (.Y(n515), 
	.A(n86));
   AND2X1 U599 (.Y(n144), 
	.B(n683), 
	.A(mem[62]));
   INVX1 U600 (.Y(n516), 
	.A(n144));
   AND2X1 U601 (.Y(n156), 
	.B(n683), 
	.A(mem[50]));
   INVX1 U602 (.Y(n517), 
	.A(n156));
   AND2X1 U603 (.Y(n106), 
	.B(FE_OFCN26_n105), 
	.A(mem[95]));
   INVX1 U604 (.Y(n518), 
	.A(n106));
   AND2X1 U605 (.Y(n119), 
	.B(FE_OFCN26_n105), 
	.A(mem[83]));
   INVX1 U606 (.Y(n519), 
	.A(n119));
   AND2X1 U607 (.Y(n213), 
	.B(n681), 
	.A(mem[5]));
   INVX1 U608 (.Y(n520), 
	.A(n213));
   AND2X1 U609 (.Y(n127), 
	.B(FE_OFCN28_n123), 
	.A(mem[76]));
   INVX1 U610 (.Y(n521), 
	.A(n127));
   AND2X1 U611 (.Y(n135), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(mem[68]));
   INVX1 U612 (.Y(n522), 
	.A(n135));
   AND2X1 U613 (.Y(n190), 
	.B(n181), 
	.A(FE_PHN72_mem_23_));
   INVX1 U614 (.Y(n523), 
	.A(n190));
   AND2X1 U615 (.Y(n171), 
	.B(n682), 
	.A(mem[38]));
   INVX1 U616 (.Y(n524), 
	.A(n171));
   AND2X1 U617 (.Y(n103), 
	.B(n684), 
	.A(mem[97]));
   INVX1 U618 (.Y(n525), 
	.A(n103));
   AND2X1 U619 (.Y(n87), 
	.B(FE_OFCN29_n55), 
	.A(mem[112]));
   INVX1 U620 (.Y(n526), 
	.A(n87));
   AND2X1 U621 (.Y(n143), 
	.B(n683), 
	.A(mem[63]));
   INVX1 U622 (.Y(n527), 
	.A(n143));
   AND2X1 U623 (.Y(n155), 
	.B(n683), 
	.A(mem[51]));
   INVX1 U624 (.Y(n528), 
	.A(n155));
   AND2X1 U625 (.Y(n107), 
	.B(FE_OFCN26_n105), 
	.A(mem[94]));
   INVX1 U626 (.Y(n529), 
	.A(n107));
   AND2X1 U627 (.Y(n120), 
	.B(FE_OFCN26_n105), 
	.A(mem[82]));
   INVX1 U628 (.Y(n530), 
	.A(n120));
   AND2X1 U629 (.Y(n212), 
	.B(n681), 
	.A(mem[6]));
   INVX1 U630 (.Y(n531), 
	.A(n212));
   AND2X1 U631 (.Y(n128), 
	.B(FE_OFCN28_n123), 
	.A(mem[75]));
   INVX1 U632 (.Y(n532), 
	.A(n128));
   AND2X2 U633 (.Y(n132), 
	.B(FE_PSN39_FE_OFCN28_n123), 
	.A(FE_PHN80_mem_71_));
   INVX1 U634 (.Y(n533), 
	.A(n132));
   AND2X2 U635 (.Y(n193), 
	.B(n181), 
	.A(FE_PHN75_mem_20_));
   INVX2 U636 (.Y(n534), 
	.A(n193));
   AND2X1 U637 (.Y(n172), 
	.B(n682), 
	.A(mem[37]));
   INVX1 U638 (.Y(n535), 
	.A(n172));
   AND2X1 U639 (.Y(n89), 
	.B(n684), 
	.A(mem[111]));
   INVX1 U640 (.Y(n536), 
	.A(n89));
   AND2X1 U641 (.Y(n102), 
	.B(n684), 
	.A(mem[98]));
   INVX1 U642 (.Y(n537), 
	.A(n102));
   AND2X1 U643 (.Y(n57), 
	.B(FE_OFCN29_n55), 
	.A(mem[126]));
   INVX1 U644 (.Y(n538), 
	.A(n57));
   AND2X2 U645 (.Y(n84), 
	.B(FE_OFCN29_n55), 
	.A(mem[115]));
   INVX1 U646 (.Y(n539), 
	.A(n84));
   AND2X1 U647 (.Y(n158), 
	.B(n683), 
	.A(mem[48]));
   INVX1 U648 (.Y(n540), 
	.A(n158));
   AND2X1 U649 (.Y(n121), 
	.B(FE_OFCN26_n105), 
	.A(mem[81]));
   INVX1 U650 (.Y(n541), 
	.A(n121));
   AND2X1 U651 (.Y(n248), 
	.B(FE_PSN47_n686), 
	.A(n685));
   INVX1 U652 (.Y(n542), 
	.A(n248));
   AND2X1 U654 (.Y(n211), 
	.B(n681), 
	.A(mem[7]));
   INVX1 U655 (.Y(n544), 
	.A(n211));
   AND2X1 U656 (.Y(n129), 
	.B(FE_OFCN28_n123), 
	.A(mem[74]));
   INVX1 U657 (.Y(n545), 
	.A(n129));
   AND2X1 U658 (.Y(n133), 
	.B(FE_OFCN28_n123), 
	.A(mem[70]));
   INVX1 U659 (.Y(n546), 
	.A(n133));
   AND2X1 U660 (.Y(n192), 
	.B(n181), 
	.A(mem[21]));
   INVX1 U661 (.Y(n547), 
	.A(n192));
   AND2X1 U662 (.Y(n173), 
	.B(n682), 
	.A(mem[36]));
   INVX1 U663 (.Y(n548), 
	.A(n173));
   AND2X1 U664 (.Y(n90), 
	.B(n684), 
	.A(mem[110]));
   INVX1 U665 (.Y(n549), 
	.A(n90));
   AND2X1 U666 (.Y(n101), 
	.B(n684), 
	.A(mem[99]));
   INVX1 U667 (.Y(n550), 
	.A(n101));
   AND2X2 U668 (.Y(n58), 
	.B(FE_PSN38_FE_OFCN29_n55), 
	.A(mem[125]));
   INVX1 U669 (.Y(n551), 
	.A(n58));
   AND2X2 U670 (.Y(n85), 
	.B(FE_PSN38_FE_OFCN29_n55), 
	.A(mem[114]));
   INVX1 U671 (.Y(n552), 
	.A(n85));
   AND2X1 U672 (.Y(n157), 
	.B(n683), 
	.A(mem[49]));
   INVX1 U673 (.Y(n553), 
	.A(n157));
   AND2X2 U674 (.Y(n122), 
	.B(FE_PSN42_FE_OFCN26_n105), 
	.A(mem[80]));
   INVX1 U675 (.Y(n554), 
	.A(n122));
   AND2X2 U676 (.Y(n220), 
	.B(n709), 
	.A(n703));
   INVX1 U677 (.Y(n555), 
	.A(n220));
   AND2X1 U678 (.Y(n160), 
	.B(n727), 
	.A(n678));
   INVX1 U679 (.Y(n556), 
	.A(n160));
   AND2X1 U680 (.Y(n180), 
	.B(n685), 
	.A(FE_PSN46_n34));
   INVX2 U681 (.Y(n557), 
	.A(n180));
   INVX8 U682 (.Y(n683), 
	.A(n558));
   INVX8 U683 (.Y(n681), 
	.A(n559));
   INVX1 U684 (.Y(n674), 
	.A(n686));
   INVX1 U685 (.Y(n675), 
	.A(FE_PSN47_n686));
   INVX1 U686 (.Y(n676), 
	.A(FE_PSN47_n686));
   INVX1 U687 (.Y(n677), 
	.A(FE_PSN47_n686));
   INVX4 U688 (.Y(n678), 
	.A(n685));
   AND2X1 U690 (.Y(n558), 
	.B(n705), 
	.A(n160));
   AND2X1 U691 (.Y(n559), 
	.B(n706), 
	.A(n237));
   INVX8 U693 (.Y(n682), 
	.A(n560));
   INVX2 U694 (.Y(n704), 
	.A(n178));
   AND2X1 U695 (.Y(n560), 
	.B(n727), 
	.A(n704));
   INVX4 U696 (.Y(n706), 
	.A(FE_OFCN20_n199));
   INVX4 U697 (.Y(n707), 
	.A(n200));
   INVX8 U698 (.Y(n684), 
	.A(n561));
   INVX2 U699 (.Y(n705), 
	.A(n159));
   INVX8 U700 (.Y(n727), 
	.A(n36));
   INVX8 U701 (.Y(n725), 
	.A(din[0]));
   INVX8 U702 (.Y(n724), 
	.A(din[1]));
   INVX8 U703 (.Y(n723), 
	.A(din[2]));
   INVX8 U704 (.Y(n722), 
	.A(din[3]));
   INVX8 U705 (.Y(n721), 
	.A(din[4]));
   INVX8 U706 (.Y(n720), 
	.A(din[5]));
   INVX8 U707 (.Y(n719), 
	.A(din[6]));
   INVX8 U708 (.Y(n718), 
	.A(din[7]));
   INVX8 U709 (.Y(n717), 
	.A(din[8]));
   INVX8 U710 (.Y(n716), 
	.A(din[9]));
   INVX8 U711 (.Y(n715), 
	.A(din[10]));
   INVX8 U712 (.Y(n714), 
	.A(din[11]));
   INVX8 U713 (.Y(n713), 
	.A(din[12]));
   INVX8 U714 (.Y(n712), 
	.A(din[13]));
   INVX8 U715 (.Y(n711), 
	.A(din[14]));
   INVX8 U716 (.Y(n710), 
	.A(din[15]));
   AND2X2 U717 (.Y(n561), 
	.B(n704), 
	.A(FE_PSN44_n36));
   INVX1 U718 (.Y(n703), 
	.A(n251));
   INVX8 U719 (.Y(n686), 
	.A(n34));
   INVX1 U720 (.Y(n702), 
	.A(FE_PHN55_FE_OFCN16_n219));
   INVX1 U721 (.Y(n64), 
	.A(n673));
   INVX1 U722 (.Y(n701), 
	.A(FE_PHN62_FE_OFCN15_n221));
   INVX1 U723 (.Y(n65), 
	.A(n672));
   INVX1 U724 (.Y(n700), 
	.A(FE_PHN64_FE_OFCN14_n222));
   INVX1 U725 (.Y(n66), 
	.A(n671));
   INVX1 U726 (.Y(n699), 
	.A(FE_PHN58_FE_OFCN13_n223));
   INVX1 U727 (.Y(n67), 
	.A(n670));
   INVX1 U728 (.Y(n698), 
	.A(FE_PHN63_FE_OFCN12_n224));
   INVX1 U729 (.Y(n68), 
	.A(n669));
   INVX1 U730 (.Y(n697), 
	.A(FE_PHN59_FE_OFCN11_n225));
   INVX1 U731 (.Y(n69), 
	.A(n668));
   INVX1 U732 (.Y(n696), 
	.A(FE_PHN61_FE_OFCN10_n226));
   INVX1 U733 (.Y(n70), 
	.A(n667));
   INVX1 U734 (.Y(n695), 
	.A(FE_PHN48_FE_OFCN9_n227));
   INVX1 U735 (.Y(n71), 
	.A(n666));
   INVX1 U736 (.Y(n694), 
	.A(FE_PHN57_FE_OFCN8_n228));
   INVX1 U737 (.Y(n72), 
	.A(n665));
   INVX1 U738 (.Y(n693), 
	.A(FE_PHN60_FE_OFCN7_n229));
   INVX1 U739 (.Y(n73), 
	.A(n664));
   INVX1 U740 (.Y(n692), 
	.A(FE_PHN53_FE_OFCN6_n230));
   INVX1 U741 (.Y(n74), 
	.A(n663));
   INVX1 U742 (.Y(n691), 
	.A(FE_PHN65_FE_OFCN5_n231));
   INVX1 U743 (.Y(n75), 
	.A(n662));
   INVX1 U744 (.Y(n690), 
	.A(FE_PHN51_FE_OFCN4_n232));
   INVX1 U745 (.Y(n76), 
	.A(n661));
   INVX1 U746 (.Y(n689), 
	.A(FE_PHN50_FE_OFCN3_n233));
   INVX1 U747 (.Y(n77), 
	.A(n660));
   INVX1 U748 (.Y(n688), 
	.A(FE_PHN52_FE_OFCN2_n234));
   INVX1 U749 (.Y(n78), 
	.A(n659));
   INVX1 U750 (.Y(n687), 
	.A(FE_PHN49_FE_OFCN1_n235));
   INVX1 U751 (.Y(n79), 
	.A(n658));
   INVX4 U752 (.Y(n685), 
	.A(n35));
   INVX8 U753 (.Y(n709), 
	.A(reset));
   INVX4 U754 (.Y(n708), 
	.A(push));
   INVX4 U755 (.Y(n726), 
	.A(empty));
   MUX2X1 U756 (.Y(n562), 
	.S(n678), 
	.B(n563), 
	.A(n564));
   MUX2X1 U757 (.Y(n565), 
	.S(n678), 
	.B(n566), 
	.A(n567));
   MUX2X1 U758 (.Y(n568), 
	.S(n678), 
	.B(n569), 
	.A(n570));
   MUX2X1 U759 (.Y(n571), 
	.S(n678), 
	.B(n572), 
	.A(n573));
   MUX2X1 U760 (.Y(n574), 
	.S(n678), 
	.B(n575), 
	.A(n576));
   MUX2X1 U761 (.Y(n577), 
	.S(n678), 
	.B(n578), 
	.A(n579));
   MUX2X1 U762 (.Y(n580), 
	.S(n678), 
	.B(n581), 
	.A(n582));
   MUX2X1 U763 (.Y(n583), 
	.S(n678), 
	.B(n584), 
	.A(n585));
   MUX2X1 U764 (.Y(n586), 
	.S(n678), 
	.B(n587), 
	.A(n588));
   MUX2X1 U765 (.Y(n589), 
	.S(n678), 
	.B(n590), 
	.A(n591));
   MUX2X1 U766 (.Y(n592), 
	.S(n678), 
	.B(n593), 
	.A(n594));
   MUX2X1 U767 (.Y(n595), 
	.S(n678), 
	.B(n596), 
	.A(n597));
   MUX2X1 U768 (.Y(n598), 
	.S(n678), 
	.B(n599), 
	.A(n600));
   MUX2X1 U769 (.Y(n601), 
	.S(n678), 
	.B(n602), 
	.A(n603));
   MUX2X1 U770 (.Y(n604), 
	.S(n678), 
	.B(n605), 
	.A(n606));
   MUX2X1 U771 (.Y(n607), 
	.S(n678), 
	.B(n608), 
	.A(n609));
   MUX2X1 U772 (.Y(n610), 
	.S(n678), 
	.B(n611), 
	.A(n612));
   MUX2X1 U773 (.Y(n613), 
	.S(n678), 
	.B(n614), 
	.A(n615));
   MUX2X1 U774 (.Y(n616), 
	.S(n678), 
	.B(n617), 
	.A(n618));
   MUX2X1 U775 (.Y(n619), 
	.S(n678), 
	.B(n620), 
	.A(n621));
   MUX2X1 U776 (.Y(n622), 
	.S(n678), 
	.B(n623), 
	.A(n624));
   MUX2X1 U777 (.Y(n625), 
	.S(n678), 
	.B(n626), 
	.A(n627));
   MUX2X1 U778 (.Y(n628), 
	.S(n678), 
	.B(n629), 
	.A(n630));
   MUX2X1 U779 (.Y(n631), 
	.S(n678), 
	.B(n632), 
	.A(n633));
   MUX2X1 U780 (.Y(n634), 
	.S(n678), 
	.B(n635), 
	.A(n636));
   MUX2X1 U781 (.Y(n637), 
	.S(n678), 
	.B(n638), 
	.A(n639));
   MUX2X1 U782 (.Y(n640), 
	.S(n678), 
	.B(n641), 
	.A(n642));
   MUX2X1 U783 (.Y(n643), 
	.S(n678), 
	.B(n644), 
	.A(n645));
   MUX2X1 U784 (.Y(n646), 
	.S(n678), 
	.B(n647), 
	.A(n648));
   MUX2X1 U785 (.Y(n649), 
	.S(n678), 
	.B(n650), 
	.A(n651));
   MUX2X1 U786 (.Y(n652), 
	.S(n678), 
	.B(n653), 
	.A(n654));
   MUX2X1 U787 (.Y(n655), 
	.S(n678), 
	.B(n656), 
	.A(n657));
   MUX2X1 U788 (.Y(n564), 
	.S(n677), 
	.B(mem[96]), 
	.A(mem[112]));
   MUX2X1 U789 (.Y(n563), 
	.S(n677), 
	.B(mem[64]), 
	.A(mem[80]));
   MUX2X1 U790 (.Y(n567), 
	.S(n677), 
	.B(mem[32]), 
	.A(mem[48]));
   MUX2X1 U791 (.Y(n566), 
	.S(n677), 
	.B(mem[0]), 
	.A(mem[16]));
   MUX2X1 U792 (.Y(n658), 
	.S(FE_PSN43_n36), 
	.B(n565), 
	.A(n562));
   MUX2X1 U793 (.Y(n570), 
	.S(n677), 
	.B(mem[97]), 
	.A(mem[113]));
   MUX2X1 U794 (.Y(n569), 
	.S(n677), 
	.B(mem[65]), 
	.A(mem[81]));
   MUX2X1 U795 (.Y(n573), 
	.S(n677), 
	.B(mem[33]), 
	.A(mem[49]));
   MUX2X1 U796 (.Y(n572), 
	.S(n677), 
	.B(mem[1]), 
	.A(mem[17]));
   MUX2X1 U797 (.Y(n659), 
	.S(FE_PSN43_n36), 
	.B(n571), 
	.A(n568));
   MUX2X1 U798 (.Y(n576), 
	.S(n677), 
	.B(mem[98]), 
	.A(mem[114]));
   MUX2X1 U799 (.Y(n575), 
	.S(n677), 
	.B(mem[66]), 
	.A(mem[82]));
   MUX2X1 U800 (.Y(n579), 
	.S(n677), 
	.B(mem[34]), 
	.A(mem[50]));
   MUX2X1 U801 (.Y(n578), 
	.S(n677), 
	.B(mem[2]), 
	.A(mem[18]));
   MUX2X1 U802 (.Y(n660), 
	.S(FE_PSN43_n36), 
	.B(n577), 
	.A(n574));
   MUX2X1 U803 (.Y(n582), 
	.S(n676), 
	.B(mem[99]), 
	.A(mem[115]));
   MUX2X1 U804 (.Y(n581), 
	.S(n676), 
	.B(mem[67]), 
	.A(mem[83]));
   MUX2X1 U805 (.Y(n585), 
	.S(n676), 
	.B(mem[35]), 
	.A(mem[51]));
   MUX2X1 U806 (.Y(n584), 
	.S(n676), 
	.B(mem[3]), 
	.A(mem[19]));
   MUX2X1 U807 (.Y(n661), 
	.S(n36), 
	.B(n583), 
	.A(n580));
   MUX2X1 U808 (.Y(n588), 
	.S(n676), 
	.B(mem[100]), 
	.A(mem[116]));
   MUX2X1 U809 (.Y(n587), 
	.S(n676), 
	.B(mem[68]), 
	.A(mem[84]));
   MUX2X1 U810 (.Y(n591), 
	.S(n676), 
	.B(mem[36]), 
	.A(mem[52]));
   MUX2X1 U811 (.Y(n590), 
	.S(n676), 
	.B(mem[4]), 
	.A(mem[20]));
   MUX2X1 U812 (.Y(n662), 
	.S(FE_PSN43_n36), 
	.B(n589), 
	.A(n586));
   MUX2X1 U813 (.Y(n594), 
	.S(n676), 
	.B(mem[101]), 
	.A(mem[117]));
   MUX2X1 U814 (.Y(n593), 
	.S(n676), 
	.B(mem[69]), 
	.A(mem[85]));
   MUX2X1 U815 (.Y(n597), 
	.S(n676), 
	.B(mem[37]), 
	.A(mem[53]));
   MUX2X1 U816 (.Y(n596), 
	.S(n676), 
	.B(mem[5]), 
	.A(mem[21]));
   MUX2X1 U817 (.Y(n663), 
	.S(FE_PSN43_n36), 
	.B(n595), 
	.A(n592));
   MUX2X1 U818 (.Y(n600), 
	.S(n675), 
	.B(mem[102]), 
	.A(mem[118]));
   MUX2X1 U819 (.Y(n599), 
	.S(n675), 
	.B(mem[70]), 
	.A(mem[86]));
   MUX2X1 U820 (.Y(n603), 
	.S(n675), 
	.B(mem[38]), 
	.A(mem[54]));
   MUX2X1 U821 (.Y(n602), 
	.S(n675), 
	.B(mem[6]), 
	.A(mem[22]));
   MUX2X1 U822 (.Y(n664), 
	.S(FE_PSN43_n36), 
	.B(n601), 
	.A(n598));
   MUX2X1 U823 (.Y(n606), 
	.S(n675), 
	.B(mem[103]), 
	.A(mem[119]));
   MUX2X1 U824 (.Y(n605), 
	.S(n675), 
	.B(mem[71]), 
	.A(mem[87]));
   MUX2X1 U825 (.Y(n609), 
	.S(n675), 
	.B(mem[39]), 
	.A(mem[55]));
   MUX2X1 U826 (.Y(n608), 
	.S(n675), 
	.B(mem[7]), 
	.A(mem[23]));
   MUX2X1 U827 (.Y(n665), 
	.S(FE_PSN43_n36), 
	.B(n607), 
	.A(n604));
   MUX2X1 U828 (.Y(n612), 
	.S(n675), 
	.B(mem[104]), 
	.A(mem[120]));
   MUX2X1 U829 (.Y(n611), 
	.S(n675), 
	.B(mem[72]), 
	.A(mem[88]));
   MUX2X1 U830 (.Y(n615), 
	.S(n675), 
	.B(mem[40]), 
	.A(mem[56]));
   MUX2X1 U831 (.Y(n614), 
	.S(n675), 
	.B(mem[8]), 
	.A(mem[24]));
   MUX2X1 U832 (.Y(n666), 
	.S(FE_PSN43_n36), 
	.B(n613), 
	.A(n610));
   MUX2X1 U833 (.Y(n618), 
	.S(n674), 
	.B(mem[105]), 
	.A(mem[121]));
   MUX2X1 U834 (.Y(n617), 
	.S(n674), 
	.B(mem[73]), 
	.A(mem[89]));
   MUX2X1 U835 (.Y(n621), 
	.S(n674), 
	.B(mem[41]), 
	.A(mem[57]));
   MUX2X1 U836 (.Y(n620), 
	.S(n674), 
	.B(mem[9]), 
	.A(mem[25]));
   MUX2X1 U837 (.Y(n667), 
	.S(FE_PSN43_n36), 
	.B(n619), 
	.A(n616));
   MUX2X1 U838 (.Y(n624), 
	.S(n674), 
	.B(mem[106]), 
	.A(mem[122]));
   MUX2X1 U839 (.Y(n623), 
	.S(n674), 
	.B(mem[74]), 
	.A(mem[90]));
   MUX2X1 U840 (.Y(n627), 
	.S(n674), 
	.B(mem[42]), 
	.A(mem[58]));
   MUX2X1 U841 (.Y(n626), 
	.S(n674), 
	.B(mem[10]), 
	.A(mem[26]));
   MUX2X1 U842 (.Y(n668), 
	.S(FE_PSN43_n36), 
	.B(n625), 
	.A(n622));
   MUX2X1 U843 (.Y(n630), 
	.S(n674), 
	.B(mem[107]), 
	.A(mem[123]));
   MUX2X1 U844 (.Y(n629), 
	.S(n674), 
	.B(mem[75]), 
	.A(mem[91]));
   MUX2X1 U845 (.Y(n633), 
	.S(n674), 
	.B(mem[43]), 
	.A(mem[59]));
   MUX2X1 U846 (.Y(n632), 
	.S(n674), 
	.B(mem[11]), 
	.A(mem[27]));
   MUX2X1 U847 (.Y(n669), 
	.S(FE_PSN43_n36), 
	.B(n631), 
	.A(n628));
   MUX2X1 U848 (.Y(n636), 
	.S(n674), 
	.B(mem[108]), 
	.A(mem[124]));
   MUX2X1 U849 (.Y(n635), 
	.S(n677), 
	.B(mem[76]), 
	.A(mem[92]));
   MUX2X1 U850 (.Y(n639), 
	.S(n676), 
	.B(mem[44]), 
	.A(mem[60]));
   MUX2X1 U851 (.Y(n638), 
	.S(n675), 
	.B(mem[12]), 
	.A(mem[28]));
   MUX2X1 U852 (.Y(n670), 
	.S(FE_PSN43_n36), 
	.B(n637), 
	.A(n634));
   MUX2X1 U853 (.Y(n642), 
	.S(n677), 
	.B(mem[109]), 
	.A(mem[125]));
   MUX2X1 U854 (.Y(n641), 
	.S(n676), 
	.B(mem[77]), 
	.A(mem[93]));
   MUX2X1 U855 (.Y(n645), 
	.S(n675), 
	.B(mem[45]), 
	.A(mem[61]));
   MUX2X1 U856 (.Y(n644), 
	.S(n674), 
	.B(mem[13]), 
	.A(mem[29]));
   MUX2X1 U857 (.Y(n671), 
	.S(FE_PSN43_n36), 
	.B(n643), 
	.A(n640));
   MUX2X1 U858 (.Y(n648), 
	.S(n676), 
	.B(mem[110]), 
	.A(mem[126]));
   MUX2X1 U859 (.Y(n647), 
	.S(n675), 
	.B(mem[78]), 
	.A(mem[94]));
   MUX2X1 U860 (.Y(n651), 
	.S(n674), 
	.B(mem[46]), 
	.A(mem[62]));
   MUX2X1 U861 (.Y(n650), 
	.S(n677), 
	.B(mem[14]), 
	.A(mem[30]));
   MUX2X1 U862 (.Y(n672), 
	.S(FE_PSN43_n36), 
	.B(n649), 
	.A(n646));
   MUX2X1 U863 (.Y(n654), 
	.S(n676), 
	.B(mem[111]), 
	.A(mem[127]));
   MUX2X1 U864 (.Y(n653), 
	.S(n677), 
	.B(mem[79]), 
	.A(mem[95]));
   MUX2X1 U865 (.Y(n657), 
	.S(n674), 
	.B(mem[47]), 
	.A(mem[63]));
   MUX2X1 U866 (.Y(n656), 
	.S(n675), 
	.B(mem[15]), 
	.A(mem[31]));
   MUX2X1 U867 (.Y(n673), 
	.S(FE_PSN43_n36), 
	.B(n655), 
	.A(n652));
endmodule


module TCAM (
	reset, 
	clk, 
	DIN, 
	EN, 
	WE, 
	match, 
	match_addr);
   input reset;
   input clk;
   input [15:0] DIN;
   input EN;
   input WE;
   output match;
   output [2:0] match_addr;

   // Internal wires
   wire FE_PHN348_last_1_;
   wire FE_PHN347_last_1_;
   wire FE_PHN346_n2877;
   wire FE_PHN345_n2851;
   wire FE_PHN344_n2851;
   wire FE_PHN343_n2877;
   wire FE_PHN342_n2889;
   wire FE_PHN341_last_1_;
   wire FE_PHN340_j_3_;
   wire FE_PHN339_n2877;
   wire FE_PHN338_n2851;
   wire FE_PHN337_n86;
   wire FE_PHN336_n2878;
   wire FE_PHN335_n2879;
   wire FE_PHN334_FE_OFCN322_n882;
   wire FE_PHN333_FE_OFCN322_n882;
   wire FE_PSN332_FE_OFCN261_n888;
   wire FE_PSN331_FE_OFCN261_n888;
   wire FE_PSN330_n960;
   wire FE_PSN329_FE_OFCN261_n888;
   wire FE_PSN328_n1003;
   wire FE_PSN327_n878;
   wire FE_PSN326_n944;
   wire FE_PSN325_n991;
   wire FE_PSN324_n926;
   wire FE_PSN323_n975;
   wire FE_OFCN322_n882;
   wire FE_OFCN321_n883;
   wire FE_OFCN320_n1021;
   wire FE_OFCN319_n1371;
   wire FE_OFCN318_n1417;
   wire FE_OFCN317_n1463;
   wire FE_OFCN316_n1334;
   wire FE_OFCN315_n1671;
   wire FE_OFCN314_n1673;
   wire FE_OFCN313_n1680;
   wire FE_OFCN312_n1607;
   wire FE_OFCN311_n1609;
   wire FE_OFCN310_n1616;
   wire FE_OFCN309_n1683;
   wire FE_OFCN308_n1531;
   wire FE_OFCN307_n1685;
   wire FE_OFCN306_n1629;
   wire FE_OFCN305_n1631;
   wire FE_OFCN304_n1638;
   wire FE_OFCN303_n1650;
   wire FE_OFCN302_n1652;
   wire FE_OFCN301_n1659;
   wire FE_OFCN300_n1565;
   wire FE_OFCN299_n1567;
   wire FE_OFCN298_n1574;
   wire FE_OFCN297_n1586;
   wire FE_OFCN296_n1588;
   wire FE_OFCN295_n1595;
   wire FE_OFCN294_n1538;
   wire FE_OFCN293_n1540;
   wire FE_OFCN292_n1547;
   wire FE_OFCN291_n1335;
   wire FE_OFCN290_n1391;
   wire FE_OFCN289_n1437;
   wire FE_OFCN288_n1485;
   wire FE_OFCN287_n1553;
   wire FE_OFCN286_n1579;
   wire FE_OFCN285_n1600;
   wire FE_OFCN284_n1688;
   wire FE_OFCN283_n1621;
   wire FE_OFCN282_n1643;
   wire FE_OFCN281_n1664;
   wire FE_OFCN280_n1697;
   wire FE_OFCN279_n2996;
   wire FE_OFCN278_n2993;
   wire FE_OFCN277_n2990;
   wire FE_OFCN276_n889;
   wire FE_OFCN275_n895;
   wire FE_OFCN268_n892;
   wire FE_OFCN267_n928;
   wire FE_OFCN266_n884;
   wire FE_OFCN263_n886;
   wire FE_OFCN261_n888;
   wire FE_OFCN255_n897;
   wire FE_OFCN251_n988;
   wire FE_OFCN250_n1005;
   wire FE_OFCN249_n1040;
   wire FE_OFCN244_n1096;
   wire FE_OFCN243_n1160;
   wire FE_OFCN242_n1129;
   wire FE_OFCN241_n1289;
   wire FE_OFCN239_n1065;
   wire FE_OFCN235_n1117;
   wire FE_OFCN233_n1150;
   wire FE_OFCN232_n1053;
   wire FE_OFCN231_n1086;
   wire FE_OFCN230_n1512;
   wire FE_OFCN229_n1368;
   wire FE_OFCN228_n1369;
   wire FE_OFCN227_n1525;
   wire FE_OFCN226_n1519;
   wire FE_OFCN225_n1667;
   wire FE_OFCN224_n1670;
   wire FE_OFCN223_n1666;
   wire FE_OFCN222_n1558;
   wire FE_OFCN221_n1561;
   wire FE_OFCN220_n1582;
   wire FE_OFCN219_n1585;
   wire FE_OFCN218_n1603;
   wire FE_OFCN217_n1606;
   wire FE_OFCN216_n1625;
   wire FE_OFCN215_n1628;
   wire FE_OFCN214_n1646;
   wire FE_OFCN213_n1649;
   wire FE_OFCN212_n1691;
   wire FE_OFCN211_n1694;
   wire FE_OFCN210_n1700;
   wire FE_OFCN209_n1703;
   wire FE_OFCN208_n1557;
   wire FE_OFCN207_n1581;
   wire FE_OFCN206_n1602;
   wire FE_OFCN205_n1624;
   wire FE_OFCN204_n1645;
   wire FE_OFCN203_n1690;
   wire FE_OFCN202_n1699;
   wire FE_OFCN201_n1034;
   wire FE_OFCN200_n1523;
   wire FE_OFCN199_n1520;
   wire FE_OFCN198_n1521;
   wire FE_OFCN197_n1031;
   wire FE_OFCN196_n1515;
   wire FE_OFCN195_n1513;
   wire FE_OFCN192_n1154;
   wire FE_OFCN191_n1058;
   wire FE_OFCN190_n1057;
   wire FE_OFCN189_n1250;
   wire FE_OFCN187_n1121;
   wire FE_OFCN186_n1122;
   wire FE_OFCN185_n1517;
   wire FE_OFCN184_n1090;
   wire FE_OFCN183_n1522;
   wire FE_OFCN179_n1526;
   wire FE_OFCN178_rank_4_;
   wire FE_OFCN177_rank_3_;
   wire FE_OFCN176_rank_5_;
   wire FE_OFCN175_n3002;
   wire FE_OFCN174_rank_10_;
   wire FE_OFCN173_rank_9_;
   wire FE_OFCN172_rank_11_;
   wire FE_OFCN171_rank_7_;
   wire FE_OFCN170_rank_6_;
   wire FE_OFCN169_rank_8_;
   wire FE_OFCN168_n3001;
   wire FE_OFCN167_rank_13_;
   wire FE_OFCN166_rank_12_;
   wire FE_OFCN165_rank_14_;
   wire FE_OFCN164_rank_23_;
   wire FE_OFCN163_rank_21_;
   wire FE_OFCN162_rank_22_;
   wire FE_OFCN140_mem_50_;
   wire FE_OFCN138_mem_52_;
   wire FE_OFCN136_mem_54_;
   wire FE_OFCN135_mem_55_;
   wire FE_OFCN134_mem_56_;
   wire FE_OFCN133_mem_57_;
   wire FE_OFCN132_mem_58_;
   wire FE_OFCN131_mem_59_;
   wire FE_OFCN130_mem_60_;
   wire FE_OFCN129_mem_61_;
   wire FE_OFCN128_mem_62_;
   wire FE_OFCN126_matchN_9_;
   wire FE_OFCN125_matchN_10_;
   wire FE_OFCN124_matchN_11_;
   wire FE_OFCN123_mem_80_;
   wire FE_OFCN122_mem_81_;
   wire FE_OFCN121_mem_82_;
   wire FE_OFCN120_mem_83_;
   wire FE_OFCN119_mem_84_;
   wire FE_OFCN118_mem_85_;
   wire FE_OFCN117_mem_86_;
   wire FE_OFCN116_mem_87_;
   wire FE_OFCN115_mem_88_;
   wire FE_OFCN114_mem_89_;
   wire FE_OFCN113_mem_90_;
   wire FE_OFCN112_mem_91_;
   wire FE_OFCN111_mem_92_;
   wire FE_OFCN110_mem_93_;
   wire FE_OFCN109_mem_94_;
   wire FE_OFCN108_mem_95_;
   wire FE_OFCN107_matchN_15_;
   wire FE_OFCN106_matchN_16_;
   wire FE_OFCN105_matchN_17_;
   wire FE_OFCN104_n2999;
   wire FE_OFCN103_m;
   wire FE_OFCN102_mem_96_;
   wire FE_OFCN101_mem_97_;
   wire FE_OFCN100_mem_98_;
   wire FE_OFCN99_mem_99_;
   wire FE_OFCN98_mem_100_;
   wire FE_OFCN97_mem_101_;
   wire FE_OFCN96_mem_102_;
   wire FE_OFCN95_mem_103_;
   wire FE_OFCN94_mem_104_;
   wire FE_OFCN93_mem_106_;
   wire FE_OFCN92_mem_107_;
   wire FE_OFCN91_mem_108_;
   wire FE_OFCN90_mem_109_;
   wire FE_OFCN89_mem_110_;
   wire FE_OFCN88_mem_111_;
   wire FE_OFCN87_matchN_18_;
   wire FE_OFCN86_matchN_19_;
   wire FE_OFCN85_matchN_20_;
   wire FE_OFCN80_mem_46_;
   wire FE_OFCN73_mem_39_;
   wire FE_OFCN71_mem_37_;
   wire FE_OFCN67_mem_33_;
   wire FE_OFCN65_matchN_14_;
   wire FE_OFCN64_matchN_13_;
   wire FE_OFCN63_matchN_12_;
   wire FE_OFCN62_mem_79_;
   wire FE_OFCN61_mem_78_;
   wire FE_OFCN60_mem_77_;
   wire FE_OFCN59_mem_76_;
   wire FE_OFCN58_mem_75_;
   wire FE_OFCN57_mem_73_;
   wire FE_OFCN56_mem_72_;
   wire FE_OFCN55_mem_71_;
   wire FE_OFCN54_mem_70_;
   wire FE_OFCN53_mem_69_;
   wire FE_OFCN52_mem_68_;
   wire FE_OFCN51_mem_67_;
   wire FE_OFCN50_mem_66_;
   wire FE_OFCN49_mem_65_;
   wire FE_OFCN48_mem_64_;
   wire FE_OFCN47_rank_16_;
   wire FE_OFCN46_rank_15_;
   wire FE_OFCN45_rank_17_;
   wire FE_OFCN44_n3000;
   wire FE_OFCN43_mem_112_;
   wire FE_OFCN42_mem_113_;
   wire FE_OFCN41_mem_114_;
   wire FE_OFCN40_mem_115_;
   wire FE_OFCN39_mem_116_;
   wire FE_OFCN38_mem_117_;
   wire FE_OFCN37_mem_118_;
   wire FE_OFCN36_mem_119_;
   wire FE_OFCN35_mem_120_;
   wire FE_OFCN34_mem_121_;
   wire FE_OFCN33_mem_122_;
   wire FE_OFCN32_mem_123_;
   wire FE_OFCN31_mem_124_;
   wire FE_OFCN30_mem_125_;
   wire FE_OFCN29_mem_126_;
   wire FE_OFCN28_mem_127_;
   wire FE_OFCN27_matchN_21_;
   wire FE_OFCN26_matchN_22_;
   wire FE_OFCN25_matchN_23_;
   wire FE_OFCN24_rank_19_;
   wire FE_OFCN23_rank_18_;
   wire FE_OFCN22_rank_20_;
   wire FE_OFCN21_mem_0_;
   wire FE_OFCN17_mem_4_;
   wire FE_OFCN5_matchN_0_;
   wire FE_OFCN4_matchN_1_;
   wire FE_OFCN3_matchN_2_;
   wire FE_OFCN2_rank_2_;
   wire FE_OFCN1_rank_1_;
   wire FE_OFCN0_rank_0_;
   wire clk__L2_N0;
   wire clk__L1_N0;
   wire n84;
   wire n85;
   wire n86;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire j_3_;
   wire n87;
   wire n88;
   wire n89;
   wire m;
   wire n250;
   wire n251;
   wire n252;
   wire n868;
   wire n870;
   wire n873;
   wire n874;
   wire n876;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n895;
   wire n897;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n919;
   wire n921;
   wire n923;
   wire n925;
   wire n926;
   wire n928;
   wire n929;
   wire n930;
   wire n932;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n948;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n964;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n979;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n995;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1005;
   wire n1007;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1021;
   wire n1023;
   wire n1025;
   wire n1027;
   wire n1028;
   wire n1030;
   wire n1031;
   wire n1033;
   wire n1034;
   wire n1036;
   wire n1037;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1049;
   wire n1051;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1057;
   wire n1058;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1069;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1090;
   wire n1092;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1113;
   wire n1115;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1121;
   wire n1122;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1133;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1154;
   wire n1156;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1178;
   wire n1180;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1186;
   wire n1187;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1198;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1219;
   wire n1221;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1242;
   wire n1244;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1250;
   wire n1251;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1262;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1283;
   wire n1285;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1317;
   wire n1319;
   wire n1321;
   wire n1323;
   wire n1325;
   wire n1327;
   wire n1329;
   wire n1331;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1342;
   wire n1345;
   wire n1348;
   wire n1350;
   wire n1352;
   wire n1354;
   wire n1356;
   wire n1358;
   wire n1360;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1395;
   wire n1396;
   wire n1398;
   wire n1400;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1409;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1441;
   wire n1442;
   wire n1444;
   wire n1446;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1455;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1490;
   wire n1492;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1501;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1517;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1531;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1538;
   wire n1540;
   wire n1542;
   wire n1545;
   wire n1547;
   wire n1548;
   wire n1550;
   wire n1553;
   wire n1554;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1565;
   wire n1567;
   wire n1569;
   wire n1572;
   wire n1574;
   wire n1575;
   wire n1577;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1588;
   wire n1590;
   wire n1593;
   wire n1595;
   wire n1596;
   wire n1598;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1609;
   wire n1611;
   wire n1614;
   wire n1616;
   wire n1617;
   wire n1619;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1631;
   wire n1633;
   wire n1636;
   wire n1638;
   wire n1639;
   wire n1641;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1652;
   wire n1654;
   wire n1657;
   wire n1659;
   wire n1660;
   wire n1662;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1673;
   wire n1675;
   wire n1678;
   wire n1680;
   wire n1681;
   wire n1683;
   wire n1685;
   wire n1686;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1708;
   wire n1716;
   wire n1781;
   wire n1844;
   wire n1890;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n238;
   wire n236;
   wire n235;
   wire n233;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2246;
   wire n2247;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2304;
   wire n2309;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2383;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2396;
   wire n2398;
   wire n2400;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2415;
   wire n2417;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2501;
   wire n2502;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2537;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2586;
   wire n2592;
   wire n2594;
   wire n2595;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2622;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2699;
   wire n2730;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2749;
   wire n2751;
   wire n2752;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire [23:0] rank;
   wire [127:0] mem;
   wire [23:0] matchN;
   wire [2:0] last;

   BUFX2 FE_PHC348_last_1_ (.Y(FE_PHN348_last_1_), 
	.A(FE_PHN347_last_1_));
   CLKBUF2 FE_PHC347_last_1_ (.Y(FE_PHN347_last_1_), 
	.A(last[1]));
   BUFX2 FE_PHC346_n2877 (.Y(FE_PHN346_n2877), 
	.A(FE_PHN339_n2877));
   BUFX2 FE_PHC345_n2851 (.Y(FE_PHN345_n2851), 
	.A(FE_PHN338_n2851));
   CLKBUF3 FE_PHC344_n2851 (.Y(FE_PHN344_n2851), 
	.A(FE_PHN345_n2851));
   CLKBUF3 FE_PHC343_n2877 (.Y(FE_PHN343_n2877), 
	.A(FE_PHN346_n2877));
   BUFX2 FE_PHC342_n2889 (.Y(FE_PHN342_n2889), 
	.A(n2889));
   CLKBUF3 FE_PHC341_last_1_ (.Y(FE_PHN341_last_1_), 
	.A(FE_PHN348_last_1_));
   CLKBUF2 FE_PHC340_j_3_ (.Y(FE_PHN340_j_3_), 
	.A(j_3_));
   BUFX2 FE_PHC339_n2877 (.Y(FE_PHN339_n2877), 
	.A(n2877));
   BUFX2 FE_PHC338_n2851 (.Y(FE_PHN338_n2851), 
	.A(n2851));
   BUFX2 FE_PHC337_n86 (.Y(FE_PHN337_n86), 
	.A(n86));
   BUFX2 FE_PHC336_n2878 (.Y(FE_PHN336_n2878), 
	.A(n2878));
   BUFX2 FE_PHC335_n2879 (.Y(n2879), 
	.A(FE_PHN335_n2879));
   BUFX2 FE_PHC334_FE_OFCN322_n882 (.Y(FE_PHN334_FE_OFCN322_n882), 
	.A(FE_PHN333_FE_OFCN322_n882));
   CLKBUF3 FE_PHC333_FE_OFCN322_n882 (.Y(FE_PHN333_FE_OFCN322_n882), 
	.A(FE_OFCN322_n882));
   BUFX2 FE_PSC332_FE_OFCN261_n888 (.Y(FE_PSN332_FE_OFCN261_n888), 
	.A(FE_OFCN261_n888));
   BUFX2 FE_PSC331_FE_OFCN261_n888 (.Y(FE_PSN331_FE_OFCN261_n888), 
	.A(FE_OFCN261_n888));
   BUFX2 FE_PSC330_n960 (.Y(FE_PSN330_n960), 
	.A(n960));
   BUFX2 FE_PSC329_FE_OFCN261_n888 (.Y(FE_PSN329_FE_OFCN261_n888), 
	.A(FE_OFCN261_n888));
   BUFX2 FE_PSC328_n1003 (.Y(FE_PSN328_n1003), 
	.A(n1003));
   BUFX2 FE_PSC327_n878 (.Y(FE_PSN327_n878), 
	.A(n878));
   BUFX2 FE_PSC326_n944 (.Y(FE_PSN326_n944), 
	.A(n944));
   BUFX2 FE_PSC325_n991 (.Y(FE_PSN325_n991), 
	.A(n991));
   BUFX2 FE_PSC324_n926 (.Y(FE_PSN324_n926), 
	.A(n926));
   BUFX2 FE_PSC323_n975 (.Y(FE_PSN323_n975), 
	.A(n975));
   BUFX2 FE_OFCC322_n882 (.Y(FE_OFCN322_n882), 
	.A(n882));
   BUFX4 FE_OFCC321_n883 (.Y(FE_OFCN321_n883), 
	.A(n883));
   BUFX4 FE_OFCC320_n1021 (.Y(FE_OFCN320_n1021), 
	.A(n1021));
   BUFX4 FE_OFCC319_n1371 (.Y(FE_OFCN319_n1371), 
	.A(n1371));
   BUFX4 FE_OFCC318_n1417 (.Y(FE_OFCN318_n1417), 
	.A(n1417));
   BUFX4 FE_OFCC317_n1463 (.Y(FE_OFCN317_n1463), 
	.A(n1463));
   BUFX2 FE_OFCC316_n1334 (.Y(FE_OFCN316_n1334), 
	.A(n1334));
   BUFX2 FE_OFCC315_n1671 (.Y(FE_OFCN315_n1671), 
	.A(n1671));
   BUFX2 FE_OFCC314_n1673 (.Y(FE_OFCN314_n1673), 
	.A(n1673));
   BUFX2 FE_OFCC313_n1680 (.Y(FE_OFCN313_n1680), 
	.A(n1680));
   BUFX4 FE_OFCC312_n1607 (.Y(FE_OFCN312_n1607), 
	.A(n1607));
   BUFX2 FE_OFCC311_n1609 (.Y(FE_OFCN311_n1609), 
	.A(n1609));
   BUFX2 FE_OFCC310_n1616 (.Y(FE_OFCN310_n1616), 
	.A(n1616));
   BUFX2 FE_OFCC309_n1683 (.Y(FE_OFCN309_n1683), 
	.A(n1683));
   BUFX2 FE_OFCC308_n1531 (.Y(FE_OFCN308_n1531), 
	.A(n1531));
   BUFX2 FE_OFCC307_n1685 (.Y(FE_OFCN307_n1685), 
	.A(n1685));
   BUFX2 FE_OFCC306_n1629 (.Y(FE_OFCN306_n1629), 
	.A(n1629));
   BUFX2 FE_OFCC305_n1631 (.Y(FE_OFCN305_n1631), 
	.A(n1631));
   BUFX2 FE_OFCC304_n1638 (.Y(FE_OFCN304_n1638), 
	.A(n1638));
   BUFX4 FE_OFCC303_n1650 (.Y(FE_OFCN303_n1650), 
	.A(n1650));
   BUFX2 FE_OFCC302_n1652 (.Y(FE_OFCN302_n1652), 
	.A(n1652));
   BUFX2 FE_OFCC301_n1659 (.Y(FE_OFCN301_n1659), 
	.A(n1659));
   BUFX2 FE_OFCC300_n1565 (.Y(FE_OFCN300_n1565), 
	.A(n1565));
   BUFX2 FE_OFCC299_n1567 (.Y(FE_OFCN299_n1567), 
	.A(n1567));
   BUFX2 FE_OFCC298_n1574 (.Y(FE_OFCN298_n1574), 
	.A(n1574));
   BUFX4 FE_OFCC297_n1586 (.Y(FE_OFCN297_n1586), 
	.A(n1586));
   BUFX2 FE_OFCC296_n1588 (.Y(FE_OFCN296_n1588), 
	.A(n1588));
   BUFX2 FE_OFCC295_n1595 (.Y(FE_OFCN295_n1595), 
	.A(n1595));
   BUFX4 FE_OFCC294_n1538 (.Y(FE_OFCN294_n1538), 
	.A(n1538));
   BUFX2 FE_OFCC293_n1540 (.Y(FE_OFCN293_n1540), 
	.A(n1540));
   BUFX2 FE_OFCC292_n1547 (.Y(FE_OFCN292_n1547), 
	.A(n1547));
   BUFX4 FE_OFCC291_n1335 (.Y(FE_OFCN291_n1335), 
	.A(n1335));
   BUFX2 FE_OFCC290_n1391 (.Y(FE_OFCN290_n1391), 
	.A(n1391));
   BUFX4 FE_OFCC289_n1437 (.Y(FE_OFCN289_n1437), 
	.A(n1437));
   BUFX4 FE_OFCC288_n1485 (.Y(FE_OFCN288_n1485), 
	.A(n1485));
   BUFX2 FE_OFCC287_n1553 (.Y(FE_OFCN287_n1553), 
	.A(n1553));
   BUFX2 FE_OFCC286_n1579 (.Y(FE_OFCN286_n1579), 
	.A(n1579));
   BUFX2 FE_OFCC285_n1600 (.Y(FE_OFCN285_n1600), 
	.A(n1600));
   BUFX2 FE_OFCC284_n1688 (.Y(FE_OFCN284_n1688), 
	.A(n1688));
   BUFX2 FE_OFCC283_n1621 (.Y(FE_OFCN283_n1621), 
	.A(n1621));
   BUFX2 FE_OFCC282_n1643 (.Y(FE_OFCN282_n1643), 
	.A(n1643));
   BUFX2 FE_OFCC281_n1664 (.Y(FE_OFCN281_n1664), 
	.A(n1664));
   BUFX2 FE_OFCC280_n1697 (.Y(FE_OFCN280_n1697), 
	.A(n1697));
   BUFX2 FE_OFCC279_n2996 (.Y(FE_OFCN279_n2996), 
	.A(n2996));
   BUFX2 FE_OFCC278_n2993 (.Y(FE_OFCN278_n2993), 
	.A(n2993));
   BUFX2 FE_OFCC277_n2990 (.Y(FE_OFCN277_n2990), 
	.A(n2990));
   BUFX2 FE_OFCC276_n889 (.Y(FE_OFCN276_n889), 
	.A(n889));
   BUFX4 FE_OFCC275_n895 (.Y(FE_OFCN275_n895), 
	.A(n895));
   BUFX4 FE_OFCC268_n892 (.Y(FE_OFCN268_n892), 
	.A(n892));
   BUFX4 FE_OFCC267_n928 (.Y(FE_OFCN267_n928), 
	.A(n928));
   BUFX2 FE_OFCC266_n884 (.Y(FE_OFCN266_n884), 
	.A(n884));
   BUFX4 FE_OFCC263_n886 (.Y(FE_OFCN263_n886), 
	.A(n886));
   BUFX4 FE_OFCC261_n888 (.Y(FE_OFCN261_n888), 
	.A(n888));
   BUFX4 FE_OFCC255_n897 (.Y(FE_OFCN255_n897), 
	.A(n897));
   BUFX2 FE_OFCC251_n988 (.Y(FE_OFCN251_n988), 
	.A(n988));
   BUFX4 FE_OFCC250_n1005 (.Y(FE_OFCN250_n1005), 
	.A(n1005));
   BUFX2 FE_OFCC249_n1040 (.Y(FE_OFCN249_n1040), 
	.A(n1040));
   BUFX2 FE_OFCC244_n1096 (.Y(FE_OFCN244_n1096), 
	.A(n1096));
   BUFX2 FE_OFCC243_n1160 (.Y(FE_OFCN243_n1160), 
	.A(n1160));
   BUFX2 FE_OFCC242_n1129 (.Y(FE_OFCN242_n1129), 
	.A(n1129));
   BUFX4 FE_OFCC241_n1289 (.Y(FE_OFCN241_n1289), 
	.A(n1289));
   BUFX2 FE_OFCC239_n1065 (.Y(FE_OFCN239_n1065), 
	.A(n1065));
   BUFX2 FE_OFCC235_n1117 (.Y(FE_OFCN235_n1117), 
	.A(n1117));
   BUFX2 FE_OFCC233_n1150 (.Y(FE_OFCN233_n1150), 
	.A(n1150));
   BUFX2 FE_OFCC232_n1053 (.Y(FE_OFCN232_n1053), 
	.A(n1053));
   BUFX2 FE_OFCC231_n1086 (.Y(FE_OFCN231_n1086), 
	.A(n1086));
   BUFX2 FE_OFCC230_n1512 (.Y(FE_OFCN230_n1512), 
	.A(n1512));
   BUFX2 FE_OFCC229_n1368 (.Y(FE_OFCN229_n1368), 
	.A(n1368));
   BUFX4 FE_OFCC228_n1369 (.Y(FE_OFCN228_n1369), 
	.A(n1369));
   BUFX2 FE_OFCC227_n1525 (.Y(FE_OFCN227_n1525), 
	.A(n1525));
   BUFX2 FE_OFCC226_n1519 (.Y(FE_OFCN226_n1519), 
	.A(n1519));
   BUFX2 FE_OFCC225_n1667 (.Y(FE_OFCN225_n1667), 
	.A(n1667));
   BUFX4 FE_OFCC224_n1670 (.Y(FE_OFCN224_n1670), 
	.A(n1670));
   BUFX2 FE_OFCC223_n1666 (.Y(FE_OFCN223_n1666), 
	.A(n1666));
   BUFX2 FE_OFCC222_n1558 (.Y(FE_OFCN222_n1558), 
	.A(n1558));
   BUFX4 FE_OFCC221_n1561 (.Y(FE_OFCN221_n1561), 
	.A(n1561));
   BUFX2 FE_OFCC220_n1582 (.Y(FE_OFCN220_n1582), 
	.A(n1582));
   BUFX2 FE_OFCC219_n1585 (.Y(FE_OFCN219_n1585), 
	.A(n1585));
   BUFX2 FE_OFCC218_n1603 (.Y(FE_OFCN218_n1603), 
	.A(n1603));
   BUFX4 FE_OFCC217_n1606 (.Y(FE_OFCN217_n1606), 
	.A(n1606));
   BUFX2 FE_OFCC216_n1625 (.Y(FE_OFCN216_n1625), 
	.A(n1625));
   BUFX2 FE_OFCC215_n1628 (.Y(FE_OFCN215_n1628), 
	.A(n1628));
   BUFX2 FE_OFCC214_n1646 (.Y(FE_OFCN214_n1646), 
	.A(n1646));
   BUFX2 FE_OFCC213_n1649 (.Y(FE_OFCN213_n1649), 
	.A(n1649));
   BUFX2 FE_OFCC212_n1691 (.Y(FE_OFCN212_n1691), 
	.A(n1691));
   BUFX4 FE_OFCC211_n1694 (.Y(FE_OFCN211_n1694), 
	.A(n1694));
   BUFX2 FE_OFCC210_n1700 (.Y(FE_OFCN210_n1700), 
	.A(n1700));
   BUFX4 FE_OFCC209_n1703 (.Y(FE_OFCN209_n1703), 
	.A(n1703));
   BUFX2 FE_OFCC208_n1557 (.Y(FE_OFCN208_n1557), 
	.A(n1557));
   BUFX2 FE_OFCC207_n1581 (.Y(FE_OFCN207_n1581), 
	.A(n1581));
   BUFX2 FE_OFCC206_n1602 (.Y(FE_OFCN206_n1602), 
	.A(n1602));
   BUFX2 FE_OFCC205_n1624 (.Y(FE_OFCN205_n1624), 
	.A(n1624));
   BUFX2 FE_OFCC204_n1645 (.Y(FE_OFCN204_n1645), 
	.A(n1645));
   BUFX2 FE_OFCC203_n1690 (.Y(FE_OFCN203_n1690), 
	.A(n1690));
   BUFX2 FE_OFCC202_n1699 (.Y(FE_OFCN202_n1699), 
	.A(n1699));
   BUFX2 FE_OFCC201_n1034 (.Y(FE_OFCN201_n1034), 
	.A(n1034));
   BUFX2 FE_OFCC200_n1523 (.Y(FE_OFCN200_n1523), 
	.A(n1523));
   BUFX2 FE_OFCC199_n1520 (.Y(FE_OFCN199_n1520), 
	.A(n1520));
   BUFX2 FE_OFCC198_n1521 (.Y(FE_OFCN198_n1521), 
	.A(n1521));
   BUFX2 FE_OFCC197_n1031 (.Y(FE_OFCN197_n1031), 
	.A(n1031));
   BUFX2 FE_OFCC196_n1515 (.Y(FE_OFCN196_n1515), 
	.A(n1515));
   BUFX2 FE_OFCC195_n1513 (.Y(FE_OFCN195_n1513), 
	.A(n1513));
   BUFX2 FE_OFCC192_n1154 (.Y(FE_OFCN192_n1154), 
	.A(n1154));
   BUFX2 FE_OFCC191_n1058 (.Y(FE_OFCN191_n1058), 
	.A(n1058));
   BUFX2 FE_OFCC190_n1057 (.Y(FE_OFCN190_n1057), 
	.A(n1057));
   BUFX4 FE_OFCC189_n1250 (.Y(FE_OFCN189_n1250), 
	.A(n1250));
   BUFX2 FE_OFCC187_n1121 (.Y(FE_OFCN187_n1121), 
	.A(n1121));
   BUFX2 FE_OFCC186_n1122 (.Y(FE_OFCN186_n1122), 
	.A(n1122));
   BUFX2 FE_OFCC185_n1517 (.Y(FE_OFCN185_n1517), 
	.A(n1517));
   BUFX2 FE_OFCC184_n1090 (.Y(FE_OFCN184_n1090), 
	.A(n1090));
   BUFX2 FE_OFCC183_n1522 (.Y(FE_OFCN183_n1522), 
	.A(n1522));
   BUFX2 FE_OFCC179_n1526 (.Y(FE_OFCN179_n1526), 
	.A(n1526));
   BUFX2 FE_OFCC178_rank_4_ (.Y(FE_OFCN178_rank_4_), 
	.A(rank[4]));
   BUFX2 FE_OFCC177_rank_3_ (.Y(FE_OFCN177_rank_3_), 
	.A(rank[3]));
   BUFX2 FE_OFCC176_rank_5_ (.Y(FE_OFCN176_rank_5_), 
	.A(rank[5]));
   BUFX2 FE_OFCC175_n3002 (.Y(FE_OFCN175_n3002), 
	.A(n3002));
   BUFX2 FE_OFCC174_rank_10_ (.Y(FE_OFCN174_rank_10_), 
	.A(rank[10]));
   BUFX2 FE_OFCC173_rank_9_ (.Y(FE_OFCN173_rank_9_), 
	.A(rank[9]));
   BUFX2 FE_OFCC172_rank_11_ (.Y(FE_OFCN172_rank_11_), 
	.A(rank[11]));
   BUFX2 FE_OFCC171_rank_7_ (.Y(FE_OFCN171_rank_7_), 
	.A(rank[7]));
   BUFX2 FE_OFCC170_rank_6_ (.Y(FE_OFCN170_rank_6_), 
	.A(rank[6]));
   BUFX2 FE_OFCC169_rank_8_ (.Y(FE_OFCN169_rank_8_), 
	.A(rank[8]));
   BUFX2 FE_OFCC168_n3001 (.Y(FE_OFCN168_n3001), 
	.A(n3001));
   BUFX2 FE_OFCC167_rank_13_ (.Y(FE_OFCN167_rank_13_), 
	.A(rank[13]));
   BUFX2 FE_OFCC166_rank_12_ (.Y(FE_OFCN166_rank_12_), 
	.A(rank[12]));
   BUFX2 FE_OFCC165_rank_14_ (.Y(FE_OFCN165_rank_14_), 
	.A(rank[14]));
   BUFX2 FE_OFCC164_rank_23_ (.Y(FE_OFCN164_rank_23_), 
	.A(rank[23]));
   BUFX2 FE_OFCC163_rank_21_ (.Y(FE_OFCN163_rank_21_), 
	.A(rank[21]));
   BUFX2 FE_OFCC162_rank_22_ (.Y(FE_OFCN162_rank_22_), 
	.A(rank[22]));
   BUFX2 FE_OFCC140_mem_50_ (.Y(FE_OFCN140_mem_50_), 
	.A(mem[50]));
   BUFX4 FE_OFCC138_mem_52_ (.Y(FE_OFCN138_mem_52_), 
	.A(mem[52]));
   BUFX2 FE_OFCC136_mem_54_ (.Y(FE_OFCN136_mem_54_), 
	.A(mem[54]));
   BUFX2 FE_OFCC135_mem_55_ (.Y(FE_OFCN135_mem_55_), 
	.A(mem[55]));
   BUFX4 FE_OFCC134_mem_56_ (.Y(FE_OFCN134_mem_56_), 
	.A(mem[56]));
   BUFX2 FE_OFCC133_mem_57_ (.Y(FE_OFCN133_mem_57_), 
	.A(mem[57]));
   BUFX2 FE_OFCC132_mem_58_ (.Y(FE_OFCN132_mem_58_), 
	.A(mem[58]));
   BUFX2 FE_OFCC131_mem_59_ (.Y(FE_OFCN131_mem_59_), 
	.A(mem[59]));
   BUFX4 FE_OFCC130_mem_60_ (.Y(FE_OFCN130_mem_60_), 
	.A(mem[60]));
   BUFX4 FE_OFCC129_mem_61_ (.Y(FE_OFCN129_mem_61_), 
	.A(mem[61]));
   BUFX4 FE_OFCC128_mem_62_ (.Y(FE_OFCN128_mem_62_), 
	.A(mem[62]));
   BUFX2 FE_OFCC126_matchN_9_ (.Y(FE_OFCN126_matchN_9_), 
	.A(matchN[9]));
   BUFX2 FE_OFCC125_matchN_10_ (.Y(FE_OFCN125_matchN_10_), 
	.A(matchN[10]));
   BUFX2 FE_OFCC124_matchN_11_ (.Y(FE_OFCN124_matchN_11_), 
	.A(matchN[11]));
   BUFX2 FE_OFCC123_mem_80_ (.Y(FE_OFCN123_mem_80_), 
	.A(mem[80]));
   BUFX2 FE_OFCC122_mem_81_ (.Y(FE_OFCN122_mem_81_), 
	.A(mem[81]));
   BUFX2 FE_OFCC121_mem_82_ (.Y(FE_OFCN121_mem_82_), 
	.A(mem[82]));
   BUFX2 FE_OFCC120_mem_83_ (.Y(FE_OFCN120_mem_83_), 
	.A(mem[83]));
   BUFX2 FE_OFCC119_mem_84_ (.Y(FE_OFCN119_mem_84_), 
	.A(mem[84]));
   BUFX2 FE_OFCC118_mem_85_ (.Y(FE_OFCN118_mem_85_), 
	.A(mem[85]));
   BUFX4 FE_OFCC117_mem_86_ (.Y(FE_OFCN117_mem_86_), 
	.A(mem[86]));
   BUFX2 FE_OFCC116_mem_87_ (.Y(FE_OFCN116_mem_87_), 
	.A(mem[87]));
   BUFX2 FE_OFCC115_mem_88_ (.Y(FE_OFCN115_mem_88_), 
	.A(mem[88]));
   BUFX2 FE_OFCC114_mem_89_ (.Y(FE_OFCN114_mem_89_), 
	.A(mem[89]));
   BUFX4 FE_OFCC113_mem_90_ (.Y(FE_OFCN113_mem_90_), 
	.A(mem[90]));
   BUFX2 FE_OFCC112_mem_91_ (.Y(FE_OFCN112_mem_91_), 
	.A(mem[91]));
   BUFX4 FE_OFCC111_mem_92_ (.Y(FE_OFCN111_mem_92_), 
	.A(mem[92]));
   BUFX2 FE_OFCC110_mem_93_ (.Y(FE_OFCN110_mem_93_), 
	.A(mem[93]));
   BUFX2 FE_OFCC109_mem_94_ (.Y(FE_OFCN109_mem_94_), 
	.A(mem[94]));
   BUFX2 FE_OFCC108_mem_95_ (.Y(FE_OFCN108_mem_95_), 
	.A(mem[95]));
   BUFX4 FE_OFCC107_matchN_15_ (.Y(FE_OFCN107_matchN_15_), 
	.A(matchN[15]));
   BUFX2 FE_OFCC106_matchN_16_ (.Y(FE_OFCN106_matchN_16_), 
	.A(matchN[16]));
   BUFX2 FE_OFCC105_matchN_17_ (.Y(FE_OFCN105_matchN_17_), 
	.A(matchN[17]));
   BUFX4 FE_OFCC104_n2999 (.Y(FE_OFCN104_n2999), 
	.A(n2999));
   BUFX2 FE_OFCC103_m (.Y(FE_OFCN103_m), 
	.A(m));
   BUFX2 FE_OFCC102_mem_96_ (.Y(FE_OFCN102_mem_96_), 
	.A(mem[96]));
   BUFX2 FE_OFCC101_mem_97_ (.Y(FE_OFCN101_mem_97_), 
	.A(mem[97]));
   BUFX2 FE_OFCC100_mem_98_ (.Y(FE_OFCN100_mem_98_), 
	.A(mem[98]));
   BUFX2 FE_OFCC99_mem_99_ (.Y(FE_OFCN99_mem_99_), 
	.A(mem[99]));
   BUFX2 FE_OFCC98_mem_100_ (.Y(FE_OFCN98_mem_100_), 
	.A(mem[100]));
   BUFX2 FE_OFCC97_mem_101_ (.Y(FE_OFCN97_mem_101_), 
	.A(mem[101]));
   BUFX2 FE_OFCC96_mem_102_ (.Y(FE_OFCN96_mem_102_), 
	.A(mem[102]));
   BUFX2 FE_OFCC95_mem_103_ (.Y(FE_OFCN95_mem_103_), 
	.A(mem[103]));
   BUFX4 FE_OFCC94_mem_104_ (.Y(FE_OFCN94_mem_104_), 
	.A(mem[104]));
   BUFX4 FE_OFCC93_mem_106_ (.Y(FE_OFCN93_mem_106_), 
	.A(mem[106]));
   BUFX2 FE_OFCC92_mem_107_ (.Y(FE_OFCN92_mem_107_), 
	.A(mem[107]));
   BUFX2 FE_OFCC91_mem_108_ (.Y(FE_OFCN91_mem_108_), 
	.A(mem[108]));
   BUFX2 FE_OFCC90_mem_109_ (.Y(FE_OFCN90_mem_109_), 
	.A(mem[109]));
   BUFX2 FE_OFCC89_mem_110_ (.Y(FE_OFCN89_mem_110_), 
	.A(mem[110]));
   BUFX2 FE_OFCC88_mem_111_ (.Y(FE_OFCN88_mem_111_), 
	.A(mem[111]));
   BUFX2 FE_OFCC87_matchN_18_ (.Y(FE_OFCN87_matchN_18_), 
	.A(matchN[18]));
   BUFX2 FE_OFCC86_matchN_19_ (.Y(FE_OFCN86_matchN_19_), 
	.A(matchN[19]));
   BUFX4 FE_OFCC85_matchN_20_ (.Y(FE_OFCN85_matchN_20_), 
	.A(matchN[20]));
   BUFX4 FE_OFCC80_mem_46_ (.Y(FE_OFCN80_mem_46_), 
	.A(mem[46]));
   BUFX2 FE_OFCC73_mem_39_ (.Y(FE_OFCN73_mem_39_), 
	.A(mem[39]));
   BUFX2 FE_OFCC71_mem_37_ (.Y(FE_OFCN71_mem_37_), 
	.A(mem[37]));
   BUFX2 FE_OFCC67_mem_33_ (.Y(FE_OFCN67_mem_33_), 
	.A(mem[33]));
   BUFX4 FE_OFCC65_matchN_14_ (.Y(FE_OFCN65_matchN_14_), 
	.A(matchN[14]));
   BUFX4 FE_OFCC64_matchN_13_ (.Y(FE_OFCN64_matchN_13_), 
	.A(matchN[13]));
   BUFX4 FE_OFCC63_matchN_12_ (.Y(FE_OFCN63_matchN_12_), 
	.A(matchN[12]));
   BUFX4 FE_OFCC62_mem_79_ (.Y(FE_OFCN62_mem_79_), 
	.A(mem[79]));
   BUFX2 FE_OFCC61_mem_78_ (.Y(FE_OFCN61_mem_78_), 
	.A(mem[78]));
   BUFX2 FE_OFCC60_mem_77_ (.Y(FE_OFCN60_mem_77_), 
	.A(mem[77]));
   BUFX2 FE_OFCC59_mem_76_ (.Y(FE_OFCN59_mem_76_), 
	.A(mem[76]));
   BUFX4 FE_OFCC58_mem_75_ (.Y(FE_OFCN58_mem_75_), 
	.A(mem[75]));
   BUFX4 FE_OFCC57_mem_73_ (.Y(FE_OFCN57_mem_73_), 
	.A(mem[73]));
   BUFX4 FE_OFCC56_mem_72_ (.Y(FE_OFCN56_mem_72_), 
	.A(mem[72]));
   BUFX4 FE_OFCC55_mem_71_ (.Y(FE_OFCN55_mem_71_), 
	.A(mem[71]));
   BUFX2 FE_OFCC54_mem_70_ (.Y(FE_OFCN54_mem_70_), 
	.A(mem[70]));
   BUFX2 FE_OFCC53_mem_69_ (.Y(FE_OFCN53_mem_69_), 
	.A(mem[69]));
   BUFX2 FE_OFCC52_mem_68_ (.Y(FE_OFCN52_mem_68_), 
	.A(mem[68]));
   BUFX2 FE_OFCC51_mem_67_ (.Y(FE_OFCN51_mem_67_), 
	.A(mem[67]));
   BUFX2 FE_OFCC50_mem_66_ (.Y(FE_OFCN50_mem_66_), 
	.A(mem[66]));
   BUFX2 FE_OFCC49_mem_65_ (.Y(FE_OFCN49_mem_65_), 
	.A(mem[65]));
   BUFX2 FE_OFCC48_mem_64_ (.Y(FE_OFCN48_mem_64_), 
	.A(mem[64]));
   BUFX4 FE_OFCC47_rank_16_ (.Y(FE_OFCN47_rank_16_), 
	.A(rank[16]));
   BUFX2 FE_OFCC46_rank_15_ (.Y(FE_OFCN46_rank_15_), 
	.A(rank[15]));
   BUFX2 FE_OFCC45_rank_17_ (.Y(FE_OFCN45_rank_17_), 
	.A(rank[17]));
   BUFX4 FE_OFCC44_n3000 (.Y(FE_OFCN44_n3000), 
	.A(n3000));
   BUFX2 FE_OFCC43_mem_112_ (.Y(FE_OFCN43_mem_112_), 
	.A(mem[112]));
   BUFX4 FE_OFCC42_mem_113_ (.Y(FE_OFCN42_mem_113_), 
	.A(mem[113]));
   BUFX2 FE_OFCC41_mem_114_ (.Y(FE_OFCN41_mem_114_), 
	.A(mem[114]));
   BUFX2 FE_OFCC40_mem_115_ (.Y(FE_OFCN40_mem_115_), 
	.A(mem[115]));
   BUFX2 FE_OFCC39_mem_116_ (.Y(FE_OFCN39_mem_116_), 
	.A(mem[116]));
   BUFX4 FE_OFCC38_mem_117_ (.Y(FE_OFCN38_mem_117_), 
	.A(mem[117]));
   BUFX2 FE_OFCC37_mem_118_ (.Y(FE_OFCN37_mem_118_), 
	.A(mem[118]));
   BUFX2 FE_OFCC36_mem_119_ (.Y(FE_OFCN36_mem_119_), 
	.A(mem[119]));
   BUFX2 FE_OFCC35_mem_120_ (.Y(FE_OFCN35_mem_120_), 
	.A(mem[120]));
   BUFX2 FE_OFCC34_mem_121_ (.Y(FE_OFCN34_mem_121_), 
	.A(mem[121]));
   BUFX2 FE_OFCC33_mem_122_ (.Y(FE_OFCN33_mem_122_), 
	.A(mem[122]));
   BUFX2 FE_OFCC32_mem_123_ (.Y(FE_OFCN32_mem_123_), 
	.A(mem[123]));
   BUFX2 FE_OFCC31_mem_124_ (.Y(FE_OFCN31_mem_124_), 
	.A(mem[124]));
   BUFX4 FE_OFCC30_mem_125_ (.Y(FE_OFCN30_mem_125_), 
	.A(mem[125]));
   BUFX2 FE_OFCC29_mem_126_ (.Y(FE_OFCN29_mem_126_), 
	.A(mem[126]));
   BUFX2 FE_OFCC28_mem_127_ (.Y(FE_OFCN28_mem_127_), 
	.A(mem[127]));
   BUFX2 FE_OFCC27_matchN_21_ (.Y(FE_OFCN27_matchN_21_), 
	.A(matchN[21]));
   BUFX2 FE_OFCC26_matchN_22_ (.Y(FE_OFCN26_matchN_22_), 
	.A(matchN[22]));
   BUFX4 FE_OFCC25_matchN_23_ (.Y(FE_OFCN25_matchN_23_), 
	.A(matchN[23]));
   BUFX2 FE_OFCC24_rank_19_ (.Y(FE_OFCN24_rank_19_), 
	.A(rank[19]));
   BUFX4 FE_OFCC23_rank_18_ (.Y(FE_OFCN23_rank_18_), 
	.A(rank[18]));
   BUFX2 FE_OFCC22_rank_20_ (.Y(FE_OFCN22_rank_20_), 
	.A(rank[20]));
   BUFX2 FE_OFCC21_mem_0_ (.Y(FE_OFCN21_mem_0_), 
	.A(mem[0]));
   BUFX2 FE_OFCC17_mem_4_ (.Y(FE_OFCN17_mem_4_), 
	.A(mem[4]));
   BUFX2 FE_OFCC5_matchN_0_ (.Y(FE_OFCN5_matchN_0_), 
	.A(matchN[0]));
   BUFX4 FE_OFCC4_matchN_1_ (.Y(FE_OFCN4_matchN_1_), 
	.A(matchN[1]));
   BUFX2 FE_OFCC3_matchN_2_ (.Y(FE_OFCN3_matchN_2_), 
	.A(matchN[2]));
   BUFX2 FE_OFCC2_rank_2_ (.Y(FE_OFCN2_rank_2_), 
	.A(rank[2]));
   BUFX2 FE_OFCC1_rank_1_ (.Y(FE_OFCN1_rank_1_), 
	.A(rank[1]));
   BUFX2 FE_OFCC0_rank_0_ (.Y(FE_OFCN0_rank_0_), 
	.A(rank[0]));
   INVX8 clk__L2_I0 (.Y(clk__L2_N0), 
	.A(clk__L1_N0));
   INVX8 clk__L1_I0 (.Y(clk__L1_N0), 
	.A(clk));
   DFFSR rank_reg_0__0_ (.S(1'b1), 
	.R(n2786), 
	.Q(rank[0]), 
	.D(n2073), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_0__1_ (.S(1'b1), 
	.R(n2779), 
	.Q(rank[1]), 
	.D(n2071), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_0__2_ (.S(1'b1), 
	.R(n2779), 
	.Q(rank[2]), 
	.D(n2070), 
	.CLK(clk__L2_N0));
   DFFPOSX1 last_reg_0_ (.Q(last[0]), 
	.D(n1899), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_0__2_ (.S(1'b1), 
	.R(n2779), 
	.Q(matchN[2]), 
	.D(n2031), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_0__1_ (.S(1'b1), 
	.R(n2779), 
	.Q(matchN[1]), 
	.D(n2032), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_0__0_ (.S(1'b1), 
	.R(n2779), 
	.Q(matchN[0]), 
	.D(n2033), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__15_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[15]), 
	.D(n2034), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__14_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[14]), 
	.D(n2035), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__13_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[13]), 
	.D(n2036), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__12_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[12]), 
	.D(n2037), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__11_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[11]), 
	.D(n2038), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__10_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[10]), 
	.D(n2039), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__9_ (.S(1'b1), 
	.R(n2779), 
	.Q(mem[9]), 
	.D(n2040), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__8_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[8]), 
	.D(n2041), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__7_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[7]), 
	.D(n2042), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__6_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[6]), 
	.D(n2043), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__5_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[5]), 
	.D(n2044), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__4_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[4]), 
	.D(n2045), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__3_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[3]), 
	.D(n2046), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__2_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[2]), 
	.D(n2047), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__1_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[1]), 
	.D(n2048), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_0__0_ (.S(1'b1), 
	.R(n2780), 
	.Q(mem[0]), 
	.D(n2049), 
	.CLK(clk__L2_N0));
   DFFPOSX1 j_reg_0_ (.Q(n84), 
	.D(n1892), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_6__2_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[20]), 
	.D(n2052), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_6__0_ (.S(1'b1), 
	.R(n2780), 
	.Q(rank[18]), 
	.D(n2054), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_6__1_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[19]), 
	.D(n2053), 
	.CLK(clk__L2_N0));
   DFFPOSX1 last_reg_2_ (.Q(last[2]), 
	.D(n1897), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_7__2_ (.S(1'b1), 
	.R(n2780), 
	.Q(matchN[23]), 
	.D(n1894), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_7__1_ (.S(1'b1), 
	.R(n2780), 
	.Q(matchN[22]), 
	.D(n1895), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_7__0_ (.S(1'b1), 
	.R(n2781), 
	.Q(matchN[21]), 
	.D(n1896), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__15_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[127]), 
	.D(n1901), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__14_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[126]), 
	.D(n1902), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__13_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[125]), 
	.D(n1903), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__12_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[124]), 
	.D(n1904), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__11_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[123]), 
	.D(n1905), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__10_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[122]), 
	.D(n1906), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__9_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[121]), 
	.D(n1907), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__8_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[120]), 
	.D(n1908), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__7_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[119]), 
	.D(n1909), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__6_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[118]), 
	.D(n1910), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__5_ (.S(1'b1), 
	.R(n2781), 
	.Q(mem[117]), 
	.D(n1911), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__4_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[116]), 
	.D(n1912), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__3_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[115]), 
	.D(n1913), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__2_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[114]), 
	.D(n1914), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__1_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[113]), 
	.D(n1915), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_7__0_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[112]), 
	.D(n1916), 
	.CLK(clk__L2_N0));
   DFFPOSX1 j_reg_2_ (.Q(n86), 
	.D(n1890), 
	.CLK(clk__L2_N0));
   DFFSR match_addr_reg_2_ (.S(1'b1), 
	.R(n2782), 
	.Q(n3000), 
	.D(n1844), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_5__2_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[17]), 
	.D(n2055), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_5__0_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[15]), 
	.D(n2057), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_5__1_ (.S(1'b1), 
	.R(n2782), 
	.Q(rank[16]), 
	.D(n2056), 
	.CLK(clk__L2_N0));
   DFFPOSX1 last_reg_1_ (.Q(last[1]), 
	.D(n1898), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__0_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[64]), 
	.D(n1973), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__1_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[65]), 
	.D(n1972), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__2_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[66]), 
	.D(n1971), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__3_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[67]), 
	.D(n1970), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__4_ (.S(1'b1), 
	.R(n2782), 
	.Q(mem[68]), 
	.D(n1969), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__5_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[69]), 
	.D(n1968), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__6_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[70]), 
	.D(n1967), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__7_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[71]), 
	.D(n1966), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__8_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[72]), 
	.D(n1965), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__9_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[73]), 
	.D(n1964), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__10_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[74]), 
	.D(n1963), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__11_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[75]), 
	.D(n1962), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__12_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[76]), 
	.D(n1961), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__13_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[77]), 
	.D(n1960), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__14_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[78]), 
	.D(n1959), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_4__15_ (.S(1'b1), 
	.R(n2783), 
	.Q(mem[79]), 
	.D(n1958), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_4__0_ (.S(1'b1), 
	.R(n2783), 
	.Q(matchN[12]), 
	.D(n1957), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_4__1_ (.S(1'b1), 
	.R(n2784), 
	.Q(matchN[13]), 
	.D(n1956), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_4__2_ (.S(1'b1), 
	.R(n2784), 
	.Q(matchN[14]), 
	.D(n1955), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__0_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[32]), 
	.D(n2011), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__1_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[33]), 
	.D(n2010), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__2_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[34]), 
	.D(n2009), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__3_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[35]), 
	.D(n2008), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__4_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[36]), 
	.D(n2007), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__5_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[37]), 
	.D(n2006), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__6_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[38]), 
	.D(n2005), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__7_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[39]), 
	.D(n2004), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__8_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[40]), 
	.D(n2003), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__9_ (.S(1'b1), 
	.R(n2784), 
	.Q(mem[41]), 
	.D(n2002), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__10_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[42]), 
	.D(n2001), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__11_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[43]), 
	.D(n2000), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__12_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[44]), 
	.D(n1999), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__13_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[45]), 
	.D(n1998), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__14_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[46]), 
	.D(n1997), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_2__15_ (.S(1'b1), 
	.R(n2785), 
	.Q(mem[47]), 
	.D(n1996), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_2__0_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[6]), 
	.D(n1995), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_2__1_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[7]), 
	.D(n1994), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_2__2_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[8]), 
	.D(n1993), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_6__2_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[20]), 
	.D(n1917), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_6__1_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[19]), 
	.D(n1918), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_6__0_ (.S(1'b1), 
	.R(n2785), 
	.Q(matchN[18]), 
	.D(n1919), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__15_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[111]), 
	.D(n1920), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__14_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[110]), 
	.D(n1921), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__13_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[109]), 
	.D(n1922), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__12_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[108]), 
	.D(n1923), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__11_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[107]), 
	.D(n1924), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__10_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[106]), 
	.D(n1925), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__9_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[105]), 
	.D(n1926), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__8_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[104]), 
	.D(n1927), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__7_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[103]), 
	.D(n1928), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__6_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[102]), 
	.D(n1929), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__5_ (.S(1'b1), 
	.R(n2786), 
	.Q(mem[101]), 
	.D(n1930), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__4_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[100]), 
	.D(n1931), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__3_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[99]), 
	.D(n1932), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__2_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[98]), 
	.D(n1933), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__1_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[97]), 
	.D(n1934), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_6__0_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[96]), 
	.D(n1935), 
	.CLK(clk__L2_N0));
   DFFSR m_reg (.S(1'b1), 
	.R(n2787), 
	.Q(m), 
	.D(n1900), 
	.CLK(clk__L2_N0));
   DFFSR match_reg (.S(1'b1), 
	.R(n2787), 
	.Q(n2999), 
	.D(n2556), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_5__2_ (.S(1'b1), 
	.R(n2787), 
	.Q(matchN[17]), 
	.D(n1936), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_5__1_ (.S(1'b1), 
	.R(n2787), 
	.Q(matchN[16]), 
	.D(n1937), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_5__0_ (.S(1'b1), 
	.R(n2787), 
	.Q(matchN[15]), 
	.D(n1938), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__15_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[95]), 
	.D(n1939), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__14_ (.S(1'b1), 
	.R(n2787), 
	.Q(mem[94]), 
	.D(n1940), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__13_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[93]), 
	.D(n1941), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__12_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[92]), 
	.D(n1942), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__11_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[91]), 
	.D(n1943), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__10_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[90]), 
	.D(n1944), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__9_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[89]), 
	.D(n1945), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__8_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[88]), 
	.D(n1946), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__7_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[87]), 
	.D(n1947), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__6_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[86]), 
	.D(n1948), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__5_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[85]), 
	.D(n1949), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__4_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[84]), 
	.D(n1950), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__3_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[83]), 
	.D(n1951), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__2_ (.S(1'b1), 
	.R(n2788), 
	.Q(mem[82]), 
	.D(n1952), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__1_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[81]), 
	.D(n1953), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_5__0_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[80]), 
	.D(n1954), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_3__2_ (.S(1'b1), 
	.R(n2789), 
	.Q(matchN[11]), 
	.D(n1974), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_3__1_ (.S(1'b1), 
	.R(n2789), 
	.Q(matchN[10]), 
	.D(n1975), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_3__0_ (.S(1'b1), 
	.R(n2789), 
	.Q(matchN[9]), 
	.D(n1976), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__15_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[63]), 
	.D(n1977), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__14_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[62]), 
	.D(n1978), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__13_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[61]), 
	.D(n1979), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__12_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[60]), 
	.D(n1980), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__11_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[59]), 
	.D(n1981), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__10_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[58]), 
	.D(n1982), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__9_ (.S(1'b1), 
	.R(n2789), 
	.Q(mem[57]), 
	.D(n1983), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__8_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[56]), 
	.D(n1984), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__7_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[55]), 
	.D(n1985), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__6_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[54]), 
	.D(n1986), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__5_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[53]), 
	.D(n1987), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__4_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[52]), 
	.D(n1988), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__3_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[51]), 
	.D(n1989), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__2_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[50]), 
	.D(n1990), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__1_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[49]), 
	.D(n1991), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_3__0_ (.S(1'b1), 
	.R(n2790), 
	.Q(mem[48]), 
	.D(n1992), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_1__2_ (.S(1'b1), 
	.R(n2790), 
	.Q(matchN[5]), 
	.D(n2012), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_1__1_ (.S(1'b1), 
	.R(n2790), 
	.Q(matchN[4]), 
	.D(n2013), 
	.CLK(clk__L2_N0));
   DFFSR matchN_reg_1__0_ (.S(1'b1), 
	.R(n2790), 
	.Q(matchN[3]), 
	.D(n2014), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__15_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[31]), 
	.D(n2015), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__14_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[30]), 
	.D(n2016), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__13_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[29]), 
	.D(n2017), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__12_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[28]), 
	.D(n2018), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__11_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[27]), 
	.D(n2019), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__10_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[26]), 
	.D(n2020), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__9_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[25]), 
	.D(n2021), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__8_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[24]), 
	.D(n2022), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__7_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[23]), 
	.D(n2023), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__6_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[22]), 
	.D(n2024), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__5_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[21]), 
	.D(n2025), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__4_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[20]), 
	.D(n2026), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__3_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[19]), 
	.D(n2027), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__2_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[18]), 
	.D(n2028), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__1_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[17]), 
	.D(n2029), 
	.CLK(clk__L2_N0));
   DFFSR mem_reg_1__0_ (.S(1'b1), 
	.R(n2796), 
	.Q(mem[16]), 
	.D(n2030), 
	.CLK(clk__L2_N0));
   DFFPOSX1 j_reg_3_ (.Q(j_3_), 
	.D(n1893), 
	.CLK(clk__L2_N0));
   DFFPOSX1 j_reg_1_ (.Q(n85), 
	.D(n2795), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_7__1_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[22]), 
	.D(n2050), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_7__0_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[21]), 
	.D(n2051), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_7__2_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[23]), 
	.D(n2072), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_4__2_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[14]), 
	.D(n2058), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_4__0_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[12]), 
	.D(n2060), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_4__1_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[13]), 
	.D(n2059), 
	.CLK(clk__L2_N0));
   DFFSR match_addr_reg_1_ (.S(1'b1), 
	.R(n2796), 
	.Q(n3001), 
	.D(n1716), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_2__2_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[8]), 
	.D(n2064), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_2__0_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[6]), 
	.D(n2066), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_2__1_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[7]), 
	.D(n2065), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_3__2_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[11]), 
	.D(n2061), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_3__0_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[9]), 
	.D(n2063), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_3__1_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[10]), 
	.D(n2062), 
	.CLK(clk__L2_N0));
   DFFSR match_addr_reg_0_ (.S(1'b1), 
	.R(n2796), 
	.Q(n3002), 
	.D(n1708), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_1__2_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[5]), 
	.D(n2067), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_1__0_ (.S(n2796), 
	.R(1'b1), 
	.Q(rank[3]), 
	.D(n2069), 
	.CLK(clk__L2_N0));
   DFFSR rank_reg_1__1_ (.S(1'b1), 
	.R(n2796), 
	.Q(rank[4]), 
	.D(n2068), 
	.CLK(clk__L2_N0));
   OAI21X1 U3 (.Y(n1708), 
	.C(n2512), 
	.B(n2871), 
	.A(n2752));
   OAI21X1 U5 (.Y(n1716), 
	.C(n2481), 
	.B(n2968), 
	.A(n2752));
   OAI21X1 U9 (.Y(n1844), 
	.C(n2447), 
	.B(n2885), 
	.A(n2752));
   OAI21X1 U12 (.Y(n1890), 
	.C(n2388), 
	.B(FE_PSN327_n878), 
	.A(n2797));
   AOI21X1 U16 (.Y(n882), 
	.C(FE_OFCN321_n883), 
	.B(n85), 
	.A(n2666));
   AOI21X1 U17 (.Y(n883), 
	.C(FE_PSN327_n878), 
	.B(n2528), 
	.A(FE_OFCN266_n884));
   NAND3X1 U18 (.Y(n884), 
	.C(FE_PSN331_FE_OFCN261_n888), 
	.B(n2502), 
	.A(FE_OFCN263_n886));
   OAI21X1 U19 (.Y(n1892), 
	.C(n2415), 
	.B(n878), 
	.A(FE_OFCN276_n889));
   AOI21X1 U22 (.Y(n889), 
	.C(n2798), 
	.B(FE_OFCN268_n892), 
	.A(n891));
   OAI21X1 U23 (.Y(n891), 
	.C(FE_OFCN263_n886), 
	.B(FE_OFCN275_n895), 
	.A(n2801));
   AOI21X1 U24 (.Y(n895), 
	.C(n2808), 
	.B(FE_OFCN255_n897), 
	.A(n2812));
   OAI21X1 U26 (.Y(n1893), 
	.C(n2434), 
	.B(n2666), 
	.A(n2844));
   OAI21X1 U29 (.Y(n901), 
	.C(n904), 
	.B(n2730), 
	.A(n902));
   NOR3X1 U30 (.Y(n902), 
	.C(n2502), 
	.B(n881), 
	.A(n2667));
   NAND3X1 U32 (.Y(n881), 
	.C(n2528), 
	.B(FE_PSN329_FE_OFCN261_n888), 
	.A(FE_OFCN263_n886));
   NAND3X1 U35 (.Y(n908), 
	.C(n911), 
	.B(n910), 
	.A(n909));
   AOI21X1 U36 (.Y(n911), 
	.C(n2501), 
	.B(FE_PHN336_n2878), 
	.A(n912));
   NAND3X1 U37 (.Y(n910), 
	.C(n917), 
	.B(n916), 
	.A(n2252));
   AOI22X1 U41 (.Y(n921), 
	.D(FE_OFCN268_n892), 
	.C(n923), 
	.B(n2309), 
	.A(n2800));
   NAND3X1 U42 (.Y(n909), 
	.C(n919), 
	.B(n2879), 
	.A(n916));
   OAI21X1 U43 (.Y(n919), 
	.C(n2244), 
	.B(FE_OFCN268_n892), 
	.A(n2929));
   OAI21X1 U47 (.Y(n912), 
	.C(FE_OFCN267_n928), 
	.B(n2928), 
	.A(FE_OFCN268_n892));
   NAND3X1 U50 (.Y(n892), 
	.C(n932), 
	.B(n930), 
	.A(n2749));
   OAI21X1 U52 (.Y(n930), 
	.C(n2928), 
	.B(n2802), 
	.A(n2803));
   AOI21X1 U55 (.Y(n928), 
	.C(n936), 
	.B(FE_OFCN105_matchN_17_), 
	.A(n2804));
   OAI21X1 U57 (.Y(n937), 
	.C(n938), 
	.B(n2929), 
	.A(FE_PSN324_n926));
   NAND3X1 U58 (.Y(n938), 
	.C(FE_OFCN87_matchN_18_), 
	.B(n2270), 
	.A(n923));
   AOI21X1 U60 (.Y(n923), 
	.C(n2247), 
	.B(n2804), 
	.A(FE_OFCN107_matchN_15_));
   OAI21X1 U63 (.Y(n926), 
	.C(n2243), 
	.B(FE_OFCN263_n886), 
	.A(n2948));
   NAND3X1 U65 (.Y(n886), 
	.C(n948), 
	.B(n946), 
	.A(n2598));
   OAI21X1 U67 (.Y(n946), 
	.C(n2947), 
	.B(n936), 
	.A(n2805));
   OAI21X1 U70 (.Y(n936), 
	.C(n952), 
	.B(n2908), 
	.A(FE_PSN329_FE_OFCN261_n888));
   OAI21X1 U72 (.Y(n953), 
	.C(n954), 
	.B(n2948), 
	.A(FE_PSN326_n944));
   NAND3X1 U73 (.Y(n954), 
	.C(FE_OFCN107_matchN_15_), 
	.B(n941), 
	.A(n2251));
   OAI21X1 U74 (.Y(n941), 
	.C(n2242), 
	.B(FE_PSN332_FE_OFCN261_n888), 
	.A(FE_OFCN63_matchN_12_));
   OAI21X1 U78 (.Y(n944), 
	.C(n2241), 
	.B(FE_PSN331_FE_OFCN261_n888), 
	.A(n2907));
   NAND3X1 U80 (.Y(n888), 
	.C(n964), 
	.B(n962), 
	.A(n2754));
   OAI21X1 U82 (.Y(n962), 
	.C(n2908), 
	.B(n2806), 
	.A(n2807));
   AOI21X1 U85 (.Y(n952), 
	.C(n967), 
	.B(FE_OFCN124_matchN_11_), 
	.A(n2808));
   OAI21X1 U87 (.Y(n968), 
	.C(n969), 
	.B(n2907), 
	.A(n960));
   NAND3X1 U88 (.Y(n969), 
	.C(FE_OFCN63_matchN_12_), 
	.B(n2269), 
	.A(n957));
   AOI21X1 U90 (.Y(n957), 
	.C(n2246), 
	.B(n2808), 
	.A(FE_OFCN126_matchN_9_));
   OAI21X1 U93 (.Y(n960), 
	.C(n2240), 
	.B(n906), 
	.A(n2955));
   NAND3X1 U95 (.Y(n906), 
	.C(n979), 
	.B(n977), 
	.A(n2586));
   OAI21X1 U97 (.Y(n977), 
	.C(n2954), 
	.B(n967), 
	.A(n2809));
   OAI21X1 U100 (.Y(n967), 
	.C(n983), 
	.B(n2927), 
	.A(FE_OFCN255_n897));
   OAI21X1 U102 (.Y(n984), 
	.C(n985), 
	.B(n2955), 
	.A(FE_PSN323_n975));
   NAND3X1 U103 (.Y(n985), 
	.C(FE_OFCN126_matchN_9_), 
	.B(n972), 
	.A(n2250));
   OAI21X1 U104 (.Y(n972), 
	.C(n2239), 
	.B(FE_OFCN255_n897), 
	.A(matchN[6]));
   OAI21X1 U107 (.Y(n975), 
	.C(n2238), 
	.B(FE_OFCN255_n897), 
	.A(n2926));
   NAND3X1 U109 (.Y(n897), 
	.C(n995), 
	.B(n993), 
	.A(n2751));
   OAI21X1 U111 (.Y(n993), 
	.C(n2927), 
	.B(n2811), 
	.A(n2810));
   AOI21X1 U114 (.Y(n983), 
	.C(n998), 
	.B(n2812), 
	.A(matchN[5]));
   OAI21X1 U116 (.Y(n999), 
	.C(n1000), 
	.B(n2926), 
	.A(FE_PSN325_n991));
   NAND3X1 U117 (.Y(n1000), 
	.C(matchN[6]), 
	.B(n2268), 
	.A(n988));
   AOI21X1 U119 (.Y(n988), 
	.C(n1002), 
	.B(n2812), 
	.A(matchN[3]));
   NOR3X1 U120 (.Y(n1002), 
	.C(n2854), 
	.B(n2812), 
	.A(n2537));
   OAI21X1 U122 (.Y(n991), 
	.C(n1007), 
	.B(FE_OFCN250_n1005), 
	.A(n2962));
   NAND3X1 U123 (.Y(n1007), 
	.C(FE_OFCN4_matchN_1_), 
	.B(FE_OFCN250_n1005), 
	.A(FE_PSN328_n1003));
   NAND3X1 U127 (.Y(n1005), 
	.C(n1011), 
	.B(n1010), 
	.A(n2592));
   OAI21X1 U128 (.Y(n1010), 
	.C(n1013), 
	.B(n2961), 
	.A(n998));
   AOI22X1 U129 (.Y(n1013), 
	.D(n1015), 
	.C(matchN[4]), 
	.B(n1014), 
	.A(matchN[3]));
   NAND3X1 U130 (.Y(n1015), 
	.C(FE_OFCN4_matchN_1_), 
	.B(n2267), 
	.A(n1003));
   OAI21X1 U132 (.Y(n1014), 
	.C(n1003), 
	.B(FE_OFCN5_matchN_0_), 
	.A(FE_OFCN4_matchN_1_));
   NAND3X1 U138 (.Y(n1018), 
	.C(n2854), 
	.B(n2852), 
	.A(n2853));
   OAI21X1 U140 (.Y(n1894), 
	.C(n2237), 
	.B(n2814), 
	.A(n1021));
   OAI21X1 U142 (.Y(n1895), 
	.C(n2236), 
	.B(n2813), 
	.A(n1021));
   OAI21X1 U144 (.Y(n1896), 
	.C(n2599), 
	.B(n2816), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U146 (.Y(n1897), 
	.C(n2235), 
	.B(FE_PHN343_n2877), 
	.A(n1028));
   OAI21X1 U149 (.Y(n1898), 
	.C(n2234), 
	.B(FE_PHN342_n2889), 
	.A(n1028));
   OAI21X1 U152 (.Y(n1899), 
	.C(n2233), 
	.B(FE_PHN344_n2851), 
	.A(n1028));
   NOR3X1 U155 (.Y(n1028), 
	.C(n904), 
	.B(reset), 
	.A(n2848));
   NOR3X1 U156 (.Y(n1900), 
	.C(n1039), 
	.B(WE), 
	.A(n2730));
   NOR3X1 U157 (.Y(n1039), 
	.C(n2420), 
	.B(n2421), 
	.A(FE_OFCN249_n1040));
   NOR3X1 U160 (.Y(n1044), 
	.C(n1047), 
	.B(n1046), 
	.A(n1045));
   XOR2X1 U161 (.Y(n1047), 
	.B(n2613), 
	.A(n2934));
   XOR2X1 U163 (.Y(n1046), 
	.B(n2495), 
	.A(n2935));
   OAI21X1 U165 (.Y(n1045), 
	.C(FE_OFCN232_n1053), 
	.B(n2930), 
	.A(DIN[15]));
   AOI22X1 U166 (.Y(n1053), 
	.D(n2938), 
	.C(n1055), 
	.B(mem[103]), 
	.A(n1054));
   OAI21X1 U167 (.Y(n1055), 
	.C(n2930), 
	.B(FE_OFCN191_n1058), 
	.A(FE_OFCN190_n1057));
   NAND3X1 U168 (.Y(n1058), 
	.C(n2945), 
	.B(n2943), 
	.A(n2944));
   NAND3X1 U169 (.Y(n1057), 
	.C(n2301), 
	.B(n2941), 
	.A(n2942));
   NOR3X1 U172 (.Y(n1043), 
	.C(n1067), 
	.B(n1066), 
	.A(FE_OFCN239_n1065));
   XOR2X1 U173 (.Y(n1067), 
	.B(n2524), 
	.A(n2936));
   XOR2X1 U175 (.Y(n1066), 
	.B(n2560), 
	.A(n2937));
   NAND3X1 U177 (.Y(n1065), 
	.C(n1074), 
	.B(n1073), 
	.A(n1072));
   XOR2X1 U178 (.Y(n1074), 
	.B(FE_OFCN90_mem_109_), 
	.A(n2437));
   XOR2X1 U180 (.Y(n1073), 
	.B(FE_OFCN89_mem_110_), 
	.A(n2485));
   XOR2X1 U182 (.Y(n1072), 
	.B(FE_OFCN91_mem_108_), 
	.A(n2518));
   NOR3X1 U185 (.Y(n1079), 
	.C(n1082), 
	.B(n1081), 
	.A(n1080));
   XNOR2X1 U186 (.Y(n1082), 
	.B(n2559), 
	.A(FE_OFCN32_mem_123_));
   XNOR2X1 U188 (.Y(n1081), 
	.B(n2461), 
	.A(FE_OFCN33_mem_122_));
   OAI21X1 U190 (.Y(n1080), 
	.C(FE_OFCN231_n1086), 
	.B(n2880), 
	.A(DIN[15]));
   AOI22X1 U191 (.Y(n1086), 
	.D(n2881), 
	.C(n1088), 
	.B(mem[119]), 
	.A(n1087));
   OAI21X1 U193 (.Y(n1088), 
	.C(n2880), 
	.B(n2884), 
	.A(FE_OFCN184_n1090));
   NOR3X1 U195 (.Y(n1092), 
	.C(FE_OFCN43_mem_112_), 
	.B(FE_OFCN41_mem_114_), 
	.A(FE_OFCN42_mem_113_));
   NAND3X1 U196 (.Y(n1090), 
	.C(n2396), 
	.B(n2882), 
	.A(n2883));
   NOR3X1 U202 (.Y(n1078), 
	.C(n1098), 
	.B(n1097), 
	.A(FE_OFCN244_n1096));
   XNOR2X1 U203 (.Y(n1098), 
	.B(n2670), 
	.A(FE_OFCN34_mem_121_));
   XNOR2X1 U205 (.Y(n1097), 
	.B(n2520), 
	.A(FE_OFCN35_mem_120_));
   NAND3X1 U207 (.Y(n1096), 
	.C(n1103), 
	.B(n1102), 
	.A(n1101));
   XOR2X1 U208 (.Y(n1103), 
	.B(FE_OFCN30_mem_125_), 
	.A(n2422));
   XOR2X1 U210 (.Y(n1102), 
	.B(FE_OFCN29_mem_126_), 
	.A(n2436));
   XOR2X1 U212 (.Y(n1101), 
	.B(FE_OFCN31_mem_124_), 
	.A(n2455));
   NOR3X1 U216 (.Y(n1108), 
	.C(n1111), 
	.B(n1110), 
	.A(n1109));
   XOR2X1 U217 (.Y(n1111), 
	.B(n2614), 
	.A(n2901));
   XOR2X1 U219 (.Y(n1110), 
	.B(n2464), 
	.A(n2900));
   OAI21X1 U221 (.Y(n1109), 
	.C(FE_OFCN235_n1117), 
	.B(n2905), 
	.A(DIN[15]));
   AOI22X1 U222 (.Y(n1117), 
	.D(n2897), 
	.C(n1119), 
	.B(FE_OFCN55_mem_71_), 
	.A(n1118));
   OAI21X1 U223 (.Y(n1119), 
	.C(n2905), 
	.B(FE_OFCN186_n1122), 
	.A(FE_OFCN187_n1121));
   NAND3X1 U224 (.Y(n1122), 
	.C(n2890), 
	.B(n2892), 
	.A(n2891));
   NAND3X1 U225 (.Y(n1121), 
	.C(n2300), 
	.B(n2894), 
	.A(n2893));
   NOR3X1 U228 (.Y(n1107), 
	.C(n1131), 
	.B(n1130), 
	.A(FE_OFCN242_n1129));
   XOR2X1 U229 (.Y(n1131), 
	.B(n2496), 
	.A(n2899));
   XOR2X1 U231 (.Y(n1130), 
	.B(n2561), 
	.A(n2898));
   NAND3X1 U233 (.Y(n1129), 
	.C(n1138), 
	.B(n1137), 
	.A(n1136));
   XOR2X1 U234 (.Y(n1138), 
	.B(FE_OFCN60_mem_77_), 
	.A(n2438));
   XOR2X1 U236 (.Y(n1137), 
	.B(FE_OFCN61_mem_78_), 
	.A(n2457));
   XOR2X1 U238 (.Y(n1136), 
	.B(FE_OFCN59_mem_76_), 
	.A(n2487));
   NOR3X1 U241 (.Y(n1143), 
	.C(n1146), 
	.B(n1145), 
	.A(n1144));
   XNOR2X1 U242 (.Y(n1146), 
	.B(n2492), 
	.A(FE_OFCN112_mem_91_));
   XNOR2X1 U244 (.Y(n1145), 
	.B(n2462), 
	.A(FE_OFCN113_mem_90_));
   OAI21X1 U246 (.Y(n1144), 
	.C(FE_OFCN233_n1150), 
	.B(n2949), 
	.A(DIN[15]));
   AOI22X1 U247 (.Y(n1150), 
	.D(n2950), 
	.C(n1152), 
	.B(FE_OFCN116_mem_87_), 
	.A(n1151));
   OAI21X1 U249 (.Y(n1152), 
	.C(n2949), 
	.B(n2953), 
	.A(FE_OFCN192_n1154));
   NOR3X1 U251 (.Y(n1156), 
	.C(mem[80]), 
	.B(mem[82]), 
	.A(FE_OFCN122_mem_81_));
   NAND3X1 U252 (.Y(n1154), 
	.C(n2398), 
	.B(n2951), 
	.A(n2952));
   NOR3X1 U258 (.Y(n1142), 
	.C(n1162), 
	.B(n1161), 
	.A(FE_OFCN243_n1160));
   XNOR2X1 U259 (.Y(n1162), 
	.B(n2671), 
	.A(FE_OFCN114_mem_89_));
   XNOR2X1 U261 (.Y(n1161), 
	.B(n2521), 
	.A(FE_OFCN115_mem_88_));
   NAND3X1 U263 (.Y(n1160), 
	.C(n1167), 
	.B(n1166), 
	.A(n1165));
   XOR2X1 U264 (.Y(n1167), 
	.B(FE_OFCN110_mem_93_), 
	.A(n2423));
   XOR2X1 U266 (.Y(n1166), 
	.B(FE_OFCN109_mem_94_), 
	.A(n2456));
   XOR2X1 U268 (.Y(n1165), 
	.B(FE_OFCN111_mem_92_), 
	.A(n2486));
   NAND3X1 U270 (.Y(n1040), 
	.C(n2299), 
	.B(n2527), 
	.A(n2468));
   NOR3X1 U273 (.Y(n1173), 
	.C(n1176), 
	.B(n1175), 
	.A(n1174));
   XOR2X1 U274 (.Y(n1176), 
	.B(n2497), 
	.A(n2858));
   XOR2X1 U276 (.Y(n1175), 
	.B(n2562), 
	.A(n2862));
   OAI21X1 U278 (.Y(n1174), 
	.C(n1182), 
	.B(n2859), 
	.A(DIN[11]));
   AOI22X1 U279 (.Y(n1182), 
	.D(n2867), 
	.C(n1184), 
	.B(mem[3]), 
	.A(n1183));
   OAI21X1 U280 (.Y(n1184), 
	.C(n2859), 
	.B(n1187), 
	.A(n1186));
   NAND3X1 U281 (.Y(n1187), 
	.C(n2870), 
	.B(n2868), 
	.A(n2869));
   NAND3X1 U282 (.Y(n1186), 
	.C(n2298), 
	.B(n2865), 
	.A(n2866));
   NOR3X1 U285 (.Y(n1172), 
	.C(n1196), 
	.B(n1195), 
	.A(n1194));
   XOR2X1 U286 (.Y(n1196), 
	.B(n2616), 
	.A(n2861));
   XOR2X1 U288 (.Y(n1195), 
	.B(n2465), 
	.A(n2860));
   NAND3X1 U290 (.Y(n1194), 
	.C(n1203), 
	.B(n1202), 
	.A(n1201));
   XOR2X1 U291 (.Y(n1203), 
	.B(mem[15]), 
	.A(n2458));
   XOR2X1 U293 (.Y(n1202), 
	.B(mem[13]), 
	.A(n2519));
   XOR2X1 U295 (.Y(n1201), 
	.B(mem[14]), 
	.A(n2488));
   NOR3X1 U298 (.Y(n1208), 
	.C(n1211), 
	.B(n1210), 
	.A(n1209));
   XNOR2X1 U299 (.Y(n1211), 
	.B(n2672), 
	.A(mem[28]));
   XNOR2X1 U301 (.Y(n1210), 
	.B(n2493), 
	.A(mem[24]));
   OAI21X1 U303 (.Y(n1209), 
	.C(n1215), 
	.B(n2963), 
	.A(DIN[11]));
   AOI22X1 U304 (.Y(n1215), 
	.D(n2966), 
	.C(n1217), 
	.B(mem[19]), 
	.A(n1216));
   OAI21X1 U306 (.Y(n1217), 
	.C(n2963), 
	.B(n2967), 
	.A(n1219));
   NOR3X1 U308 (.Y(n1221), 
	.C(mem[16]), 
	.B(mem[18]), 
	.A(mem[17]));
   NAND3X1 U309 (.Y(n1219), 
	.C(n2417), 
	.B(n2964), 
	.A(n2965));
   NOR3X1 U315 (.Y(n1207), 
	.C(n1227), 
	.B(n1226), 
	.A(n1225));
   XNOR2X1 U316 (.Y(n1227), 
	.B(n2523), 
	.A(mem[25]));
   XNOR2X1 U318 (.Y(n1226), 
	.B(n2463), 
	.A(mem[26]));
   NAND3X1 U320 (.Y(n1225), 
	.C(n1232), 
	.B(n1231), 
	.A(n1230));
   XOR2X1 U321 (.Y(n1232), 
	.B(mem[31]), 
	.A(n2439));
   XOR2X1 U323 (.Y(n1231), 
	.B(mem[29]), 
	.A(n2459));
   XOR2X1 U325 (.Y(n1230), 
	.B(mem[30]), 
	.A(n2489));
   NOR3X1 U328 (.Y(n1237), 
	.C(n1240), 
	.B(n1239), 
	.A(n1238));
   XOR2X1 U329 (.Y(n1240), 
	.B(n2615), 
	.A(n2920));
   XOR2X1 U331 (.Y(n1239), 
	.B(n2466), 
	.A(n2919));
   OAI21X1 U333 (.Y(n1238), 
	.C(n1246), 
	.B(n2924), 
	.A(DIN[15]));
   AOI22X1 U334 (.Y(n1246), 
	.D(n2916), 
	.C(n1248), 
	.B(FE_OFCN73_mem_39_), 
	.A(n1247));
   OAI21X1 U335 (.Y(n1248), 
	.C(n2924), 
	.B(n1251), 
	.A(FE_OFCN189_n1250));
   NAND3X1 U336 (.Y(n1251), 
	.C(n2909), 
	.B(n2911), 
	.A(n2910));
   NAND3X1 U337 (.Y(n1250), 
	.C(n2297), 
	.B(n2913), 
	.A(n2912));
   NOR3X1 U340 (.Y(n1236), 
	.C(n1260), 
	.B(n1259), 
	.A(n1258));
   XOR2X1 U341 (.Y(n1260), 
	.B(n2498), 
	.A(n2918));
   XOR2X1 U343 (.Y(n1259), 
	.B(n2563), 
	.A(n2917));
   NAND3X1 U345 (.Y(n1258), 
	.C(n1267), 
	.B(n1266), 
	.A(n1265));
   XOR2X1 U346 (.Y(n1267), 
	.B(mem[45]), 
	.A(n2441));
   XOR2X1 U348 (.Y(n1266), 
	.B(FE_OFCN80_mem_46_), 
	.A(n2460));
   XOR2X1 U350 (.Y(n1265), 
	.B(mem[44]), 
	.A(n2491));
   NOR3X1 U353 (.Y(n1272), 
	.C(n1275), 
	.B(n1274), 
	.A(n1273));
   XNOR2X1 U354 (.Y(n1275), 
	.B(n2494), 
	.A(FE_OFCN131_mem_59_));
   XNOR2X1 U356 (.Y(n1274), 
	.B(n2442), 
	.A(FE_OFCN132_mem_58_));
   OAI21X1 U358 (.Y(n1273), 
	.C(n1279), 
	.B(n2956), 
	.A(DIN[15]));
   AOI22X1 U359 (.Y(n1279), 
	.D(n2957), 
	.C(n1281), 
	.B(FE_OFCN135_mem_55_), 
	.A(n1280));
   OAI21X1 U361 (.Y(n1281), 
	.C(n2956), 
	.B(n2960), 
	.A(n1283));
   NOR3X1 U363 (.Y(n1285), 
	.C(mem[48]), 
	.B(mem[50]), 
	.A(mem[49]));
   NAND3X1 U364 (.Y(n1283), 
	.C(n2400), 
	.B(n2958), 
	.A(n2959));
   NOR3X1 U370 (.Y(n1271), 
	.C(n1291), 
	.B(n1290), 
	.A(FE_OFCN241_n1289));
   XNOR2X1 U371 (.Y(n1291), 
	.B(n2673), 
	.A(FE_OFCN133_mem_57_));
   XNOR2X1 U373 (.Y(n1290), 
	.B(n2522), 
	.A(FE_OFCN134_mem_56_));
   NAND3X1 U375 (.Y(n1289), 
	.C(n1296), 
	.B(n1295), 
	.A(n1294));
   XOR2X1 U376 (.Y(n1296), 
	.B(FE_OFCN129_mem_61_), 
	.A(n2424));
   XOR2X1 U378 (.Y(n1295), 
	.B(FE_OFCN128_mem_62_), 
	.A(n2440));
   XOR2X1 U380 (.Y(n1294), 
	.B(FE_OFCN130_mem_60_), 
	.A(n2490));
   OAI21X1 U382 (.Y(n1901), 
	.C(n2232), 
	.B(n2743), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U384 (.Y(n1902), 
	.C(n2231), 
	.B(n2745), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U386 (.Y(n1903), 
	.C(n2445), 
	.B(n2746), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U388 (.Y(n1904), 
	.C(n2230), 
	.B(n2744), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U390 (.Y(n1905), 
	.C(n2229), 
	.B(n2739), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U392 (.Y(n1906), 
	.C(n2387), 
	.B(n2740), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U394 (.Y(n1907), 
	.C(n2228), 
	.B(n2741), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U396 (.Y(n1908), 
	.C(n2227), 
	.B(n2742), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U398 (.Y(n1909), 
	.C(n2473), 
	.B(n2817), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U400 (.Y(n1910), 
	.C(n2545), 
	.B(n2819), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U402 (.Y(n1911), 
	.C(n2505), 
	.B(n2820), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U404 (.Y(n1912), 
	.C(n2226), 
	.B(n2821), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U406 (.Y(n1913), 
	.C(n2225), 
	.B(n2822), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U408 (.Y(n1914), 
	.C(n2407), 
	.B(n2824), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U410 (.Y(n1915), 
	.C(n2427), 
	.B(n2825), 
	.A(FE_OFCN320_n1021));
   OAI21X1 U412 (.Y(n1916), 
	.C(n2446), 
	.B(n2826), 
	.A(FE_OFCN320_n1021));
   NAND3X1 U414 (.Y(n1021), 
	.C(FE_OFCN316_n1334), 
	.B(n2847), 
	.A(n2846));
   OAI21X1 U415 (.Y(n1917), 
	.C(n2224), 
	.B(n2928), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U418 (.Y(n1918), 
	.C(n2223), 
	.B(n2929), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U421 (.Y(n1919), 
	.C(n2669), 
	.B(n2309), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U424 (.Y(n1920), 
	.C(n2222), 
	.B(n2930), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U427 (.Y(n1921), 
	.C(n2517), 
	.B(n2931), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U430 (.Y(n1922), 
	.C(n2554), 
	.B(n2932), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U433 (.Y(n1923), 
	.C(n2608), 
	.B(n2933), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U436 (.Y(n1924), 
	.C(n2221), 
	.B(n2934), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U439 (.Y(n1925), 
	.C(n2220), 
	.B(n2935), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U442 (.Y(n1926), 
	.C(n2219), 
	.B(n2936), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U445 (.Y(n1927), 
	.C(n2218), 
	.B(n2937), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U448 (.Y(n1928), 
	.C(n2391), 
	.B(n2938), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U451 (.Y(n1929), 
	.C(n2555), 
	.B(n2939), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U454 (.Y(n1930), 
	.C(n2609), 
	.B(n2940), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U457 (.Y(n1931), 
	.C(n2410), 
	.B(n2941), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U460 (.Y(n1932), 
	.C(n2430), 
	.B(n2942), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U463 (.Y(n1933), 
	.C(n2450), 
	.B(n2943), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U466 (.Y(n1934), 
	.C(n2476), 
	.B(n2944), 
	.A(FE_OFCN291_n1335));
   OAI21X1 U469 (.Y(n1935), 
	.C(n2506), 
	.B(n2945), 
	.A(FE_OFCN291_n1335));
   NOR3X1 U472 (.Y(n1335), 
	.C(n2594), 
	.B(FE_OFCN228_n1369), 
	.A(FE_OFCN229_n1368));
   OAI21X1 U473 (.Y(n1936), 
	.C(n2217), 
	.B(n1371), 
	.A(n2814));
   OAI21X1 U475 (.Y(n1937), 
	.C(n2216), 
	.B(n1371), 
	.A(n2813));
   OAI21X1 U477 (.Y(n1938), 
	.C(n2215), 
	.B(n1371), 
	.A(n2816));
   OAI21X1 U479 (.Y(n1939), 
	.C(n2214), 
	.B(FE_OFCN319_n1371), 
	.A(n2743));
   OAI21X1 U481 (.Y(n1940), 
	.C(n2213), 
	.B(FE_OFCN319_n1371), 
	.A(n2745));
   OAI21X1 U483 (.Y(n1941), 
	.C(n2507), 
	.B(FE_OFCN319_n1371), 
	.A(n2746));
   OAI21X1 U485 (.Y(n1942), 
	.C(n2212), 
	.B(FE_OFCN319_n1371), 
	.A(n2744));
   OAI21X1 U487 (.Y(n1943), 
	.C(n2211), 
	.B(FE_OFCN319_n1371), 
	.A(n2739));
   OAI21X1 U489 (.Y(n1944), 
	.C(n2411), 
	.B(FE_OFCN319_n1371), 
	.A(n2740));
   OAI21X1 U491 (.Y(n1945), 
	.C(n2392), 
	.B(n1371), 
	.A(n2741));
   OAI21X1 U493 (.Y(n1946), 
	.C(n2210), 
	.B(n1371), 
	.A(n2742));
   OAI21X1 U495 (.Y(n1947), 
	.C(n2600), 
	.B(FE_OFCN319_n1371), 
	.A(n2817));
   OAI21X1 U497 (.Y(n1948), 
	.C(n2431), 
	.B(FE_OFCN319_n1371), 
	.A(n2819));
   OAI21X1 U499 (.Y(n1949), 
	.C(n2546), 
	.B(FE_OFCN319_n1371), 
	.A(n2820));
   OAI21X1 U501 (.Y(n1950), 
	.C(n2209), 
	.B(FE_OFCN319_n1371), 
	.A(n2821));
   OAI21X1 U503 (.Y(n1951), 
	.C(n2208), 
	.B(FE_OFCN319_n1371), 
	.A(n2822));
   OAI21X1 U505 (.Y(n1952), 
	.C(n2508), 
	.B(FE_OFCN319_n1371), 
	.A(n2824));
   OAI21X1 U507 (.Y(n1953), 
	.C(n2451), 
	.B(FE_OFCN319_n1371), 
	.A(n2825));
   OAI21X1 U509 (.Y(n1954), 
	.C(n2477), 
	.B(FE_OFCN319_n1371), 
	.A(n2826));
   NAND3X1 U511 (.Y(n1371), 
	.C(FE_OFCN228_n1369), 
	.B(n2846), 
	.A(FE_OFCN316_n1334));
   OAI21X1 U512 (.Y(n1955), 
	.C(n2428), 
	.B(n2908), 
	.A(n1391));
   OAI21X1 U515 (.Y(n1956), 
	.C(n2408), 
	.B(n2907), 
	.A(n1391));
   OAI21X1 U518 (.Y(n1957), 
	.C(n2514), 
	.B(n2906), 
	.A(n1391));
   OAI21X1 U521 (.Y(n1958), 
	.C(n2389), 
	.B(n2905), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U524 (.Y(n1959), 
	.C(n2552), 
	.B(n2904), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U527 (.Y(n1960), 
	.C(n2483), 
	.B(n2903), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U530 (.Y(n1961), 
	.C(n2454), 
	.B(n2902), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U533 (.Y(n1962), 
	.C(n2448), 
	.B(n2901), 
	.A(n1391));
   OAI21X1 U536 (.Y(n1963), 
	.C(n2207), 
	.B(n2900), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U539 (.Y(n1964), 
	.C(n2206), 
	.B(n2899), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U542 (.Y(n1965), 
	.C(n2205), 
	.B(n2898), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U545 (.Y(n1966), 
	.C(n2204), 
	.B(n2897), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U548 (.Y(n1967), 
	.C(n2551), 
	.B(n2896), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U551 (.Y(n1968), 
	.C(n2605), 
	.B(n2895), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U554 (.Y(n1969), 
	.C(n2474), 
	.B(n2894), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U557 (.Y(n1970), 
	.C(n2203), 
	.B(n2893), 
	.A(FE_OFCN290_n1391));
   OAI21X1 U560 (.Y(n1971), 
	.C(n2202), 
	.B(n2892), 
	.A(n1391));
   OAI21X1 U563 (.Y(n1972), 
	.C(n2201), 
	.B(n2891), 
	.A(n1391));
   OAI21X1 U566 (.Y(n1973), 
	.C(n2200), 
	.B(n2890), 
	.A(FE_OFCN290_n1391));
   NOR3X1 U569 (.Y(n1391), 
	.C(n2847), 
	.B(FE_OFCN229_n1368), 
	.A(n2594));
   OAI21X1 U570 (.Y(n1974), 
	.C(n2199), 
	.B(n1417), 
	.A(n2814));
   OAI21X1 U572 (.Y(n1975), 
	.C(n2198), 
	.B(n1417), 
	.A(n2813));
   OAI21X1 U574 (.Y(n1976), 
	.C(n2197), 
	.B(n1417), 
	.A(n2816));
   OAI21X1 U576 (.Y(n1977), 
	.C(n2196), 
	.B(FE_OFCN318_n1417), 
	.A(n2743));
   OAI21X1 U578 (.Y(n1978), 
	.C(n2195), 
	.B(FE_OFCN318_n1417), 
	.A(n2745));
   OAI21X1 U580 (.Y(n1979), 
	.C(n2478), 
	.B(FE_OFCN318_n1417), 
	.A(n2746));
   OAI21X1 U582 (.Y(n1980), 
	.C(n2194), 
	.B(FE_OFCN318_n1417), 
	.A(n2744));
   OAI21X1 U584 (.Y(n1981), 
	.C(n2193), 
	.B(FE_OFCN318_n1417), 
	.A(n2739));
   OAI21X1 U586 (.Y(n1982), 
	.C(n2192), 
	.B(FE_OFCN318_n1417), 
	.A(n2740));
   OAI21X1 U588 (.Y(n1983), 
	.C(n2412), 
	.B(n1417), 
	.A(n2741));
   OAI21X1 U590 (.Y(n1984), 
	.C(n2393), 
	.B(n1417), 
	.A(n2742));
   OAI21X1 U592 (.Y(n1985), 
	.C(n2432), 
	.B(FE_OFCN318_n1417), 
	.A(n2817));
   OAI21X1 U594 (.Y(n1986), 
	.C(n2452), 
	.B(FE_OFCN318_n1417), 
	.A(n2819));
   OAI21X1 U596 (.Y(n1987), 
	.C(n2601), 
	.B(FE_OFCN318_n1417), 
	.A(n2820));
   OAI21X1 U598 (.Y(n1988), 
	.C(n2191), 
	.B(FE_OFCN318_n1417), 
	.A(n2821));
   OAI21X1 U600 (.Y(n1989), 
	.C(n2190), 
	.B(FE_OFCN318_n1417), 
	.A(n2822));
   OAI21X1 U602 (.Y(n1990), 
	.C(n2479), 
	.B(FE_OFCN318_n1417), 
	.A(n2824));
   OAI21X1 U604 (.Y(n1991), 
	.C(n2509), 
	.B(n1417), 
	.A(n2825));
   OAI21X1 U606 (.Y(n1992), 
	.C(n2547), 
	.B(FE_OFCN318_n1417), 
	.A(n2826));
   NAND3X1 U608 (.Y(n1417), 
	.C(FE_OFCN229_n1368), 
	.B(n2847), 
	.A(FE_OFCN316_n1334));
   OAI21X1 U609 (.Y(n1993), 
	.C(n2449), 
	.B(n2927), 
	.A(n1437));
   OAI21X1 U612 (.Y(n1994), 
	.C(n2668), 
	.B(n2926), 
	.A(n1437));
   OAI21X1 U615 (.Y(n1995), 
	.C(n2553), 
	.B(n2925), 
	.A(n1437));
   OAI21X1 U618 (.Y(n1996), 
	.C(n2429), 
	.B(n2924), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U621 (.Y(n1997), 
	.C(n2607), 
	.B(n2923), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U624 (.Y(n1998), 
	.C(n2516), 
	.B(n2922), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U627 (.Y(n1999), 
	.C(n2484), 
	.B(n2921), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U630 (.Y(n2000), 
	.C(n2475), 
	.B(n2920), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U633 (.Y(n2001), 
	.C(n2409), 
	.B(n2919), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U636 (.Y(n2002), 
	.C(n2390), 
	.B(n2918), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U639 (.Y(n2003), 
	.C(n2189), 
	.B(n2917), 
	.A(n1437));
   OAI21X1 U642 (.Y(n2004), 
	.C(n2188), 
	.B(n2916), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U645 (.Y(n2005), 
	.C(n2515), 
	.B(n2915), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U648 (.Y(n2006), 
	.C(n2606), 
	.B(n2914), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U651 (.Y(n2007), 
	.C(n2187), 
	.B(n2913), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U654 (.Y(n2008), 
	.C(n2186), 
	.B(n2912), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U657 (.Y(n2009), 
	.C(n2185), 
	.B(n2911), 
	.A(FE_OFCN289_n1437));
   OAI21X1 U660 (.Y(n2010), 
	.C(n2184), 
	.B(n2910), 
	.A(n1437));
   OAI21X1 U663 (.Y(n2011), 
	.C(n2183), 
	.B(n2909), 
	.A(FE_OFCN289_n1437));
   NOR3X1 U666 (.Y(n1437), 
	.C(n2846), 
	.B(FE_OFCN228_n1369), 
	.A(n2594));
   OAI21X1 U667 (.Y(n2012), 
	.C(n2182), 
	.B(n1463), 
	.A(n2814));
   OAI21X1 U670 (.Y(n2013), 
	.C(n2181), 
	.B(n1463), 
	.A(n2813));
   OAI21X1 U673 (.Y(n2014), 
	.C(n2180), 
	.B(n1463), 
	.A(n2816));
   OAI21X1 U676 (.Y(n2015), 
	.C(n2179), 
	.B(FE_OFCN317_n1463), 
	.A(n2743));
   OAI21X1 U678 (.Y(n2016), 
	.C(n2510), 
	.B(FE_OFCN317_n1463), 
	.A(n2745));
   OAI21X1 U680 (.Y(n2017), 
	.C(n2548), 
	.B(FE_OFCN317_n1463), 
	.A(n2746));
   OAI21X1 U682 (.Y(n2018), 
	.C(n2178), 
	.B(FE_OFCN317_n1463), 
	.A(n2744));
   OAI21X1 U684 (.Y(n2019), 
	.C(n2177), 
	.B(FE_OFCN317_n1463), 
	.A(n2739));
   OAI21X1 U686 (.Y(n2020), 
	.C(n2176), 
	.B(FE_OFCN317_n1463), 
	.A(n2740));
   OAI21X1 U688 (.Y(n2021), 
	.C(n2175), 
	.B(FE_OFCN317_n1463), 
	.A(n2741));
   OAI21X1 U690 (.Y(n2022), 
	.C(n2413), 
	.B(FE_OFCN317_n1463), 
	.A(n2742));
   OAI21X1 U692 (.Y(n2023), 
	.C(n2174), 
	.B(FE_OFCN317_n1463), 
	.A(n2817));
   OAI21X1 U695 (.Y(n2024), 
	.C(n2394), 
	.B(FE_OFCN317_n1463), 
	.A(n2819));
   OAI21X1 U698 (.Y(n2025), 
	.C(n2433), 
	.B(FE_OFCN317_n1463), 
	.A(n2820));
   OAI21X1 U701 (.Y(n2026), 
	.C(n2453), 
	.B(FE_OFCN317_n1463), 
	.A(n2821));
   OAI21X1 U704 (.Y(n2027), 
	.C(n2511), 
	.B(n1463), 
	.A(n2822));
   OAI21X1 U707 (.Y(n2028), 
	.C(n2549), 
	.B(n1463), 
	.A(n2824));
   OAI21X1 U710 (.Y(n2029), 
	.C(n2480), 
	.B(n1463), 
	.A(n2825));
   OAI21X1 U713 (.Y(n2030), 
	.C(n2602), 
	.B(n1463), 
	.A(n2826));
   NAND3X1 U715 (.Y(n1463), 
	.C(n1368), 
	.B(FE_OFCN316_n1334), 
	.A(FE_OFCN228_n1369));
   AOI21X1 U716 (.Y(n1334), 
	.C(n904), 
	.B(n2873), 
	.A(n2469));
   OAI21X1 U718 (.Y(n2031), 
	.C(n2173), 
	.B(n2852), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U721 (.Y(n2032), 
	.C(n2172), 
	.B(n2853), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U724 (.Y(n2033), 
	.C(n2171), 
	.B(n2854), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U727 (.Y(n2034), 
	.C(n2513), 
	.B(n2855), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U732 (.Y(n2035), 
	.C(n2482), 
	.B(n2856), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U737 (.Y(n2036), 
	.C(n2603), 
	.B(n2857), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U742 (.Y(n2037), 
	.C(n2425), 
	.B(n2858), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U747 (.Y(n2038), 
	.C(n2170), 
	.B(n2859), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U752 (.Y(n2039), 
	.C(n2169), 
	.B(n2860), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U757 (.Y(n2040), 
	.C(n2168), 
	.B(n2861), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U762 (.Y(n2041), 
	.C(n2167), 
	.B(n2862), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U767 (.Y(n2042), 
	.C(n2550), 
	.B(n2863), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U770 (.Y(n2043), 
	.C(n2604), 
	.B(n2864), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U773 (.Y(n2044), 
	.C(n2166), 
	.B(n2865), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U776 (.Y(n2045), 
	.C(n2386), 
	.B(n2866), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U779 (.Y(n2046), 
	.C(n2406), 
	.B(n2867), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U782 (.Y(n2047), 
	.C(n2426), 
	.B(n2868), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U785 (.Y(n2048), 
	.C(n2444), 
	.B(n2869), 
	.A(FE_OFCN288_n1485));
   OAI21X1 U788 (.Y(n2049), 
	.C(n2472), 
	.B(n2870), 
	.A(FE_OFCN288_n1485));
   NOR3X1 U791 (.Y(n1485), 
	.C(n2846), 
	.B(n2594), 
	.A(n2847));
   AOI21X1 U793 (.Y(n1368), 
	.C(FE_OFCN197_n1031), 
	.B(last[2]), 
	.A(n2848));
   OAI21X1 U798 (.Y(n1037), 
	.C(FE_OFCN195_n1513), 
	.B(FE_OFCN230_n1512), 
	.A(n2874));
   AOI21X1 U799 (.Y(n1512), 
	.C(n2383), 
	.B(FE_OFCN196_n1515), 
	.A(n1514));
   OAI21X1 U801 (.Y(n1514), 
	.C(FE_OFCN199_n1520), 
	.B(FE_OFCN226_n1519), 
	.A(n2304));
   AOI21X1 U805 (.Y(n1369), 
	.C(FE_OFCN201_n1034), 
	.B(last[1]), 
	.A(n2848));
   NAND3X1 U806 (.Y(n1034), 
	.C(FE_OFCN200_n1523), 
	.B(FE_OFCN195_n1513), 
	.A(FE_OFCN183_n1522));
   NAND3X1 U807 (.Y(n1523), 
	.C(n2351), 
	.B(FE_OFCN185_n1517), 
	.A(FE_OFCN196_n1515));
   NAND3X1 U809 (.Y(n1525), 
	.C(n2296), 
	.B(FE_OFCN226_n1519), 
	.A(FE_OFCN179_n1526));
   NAND3X1 U812 (.Y(n1520), 
	.C(FE_OFCN172_rank_11_), 
	.B(rank[9]), 
	.A(rank[10]));
   NAND3X1 U813 (.Y(n1521), 
	.C(FE_OFCN169_rank_8_), 
	.B(rank[6]), 
	.A(rank[7]));
   NAND3X1 U814 (.Y(n1031), 
	.C(n1528), 
	.B(FE_OFCN185_n1517), 
	.A(FE_OFCN196_n1515));
   NAND3X1 U816 (.Y(n1513), 
	.C(FE_OFCN164_rank_23_), 
	.B(rank[21]), 
	.A(FE_OFCN162_rank_22_));
   NAND3X1 U817 (.Y(n1522), 
	.C(FE_OFCN22_rank_20_), 
	.B(FE_OFCN23_rank_18_), 
	.A(rank[19]));
   NAND3X1 U818 (.Y(n1517), 
	.C(FE_OFCN45_rank_17_), 
	.B(FE_OFCN46_rank_15_), 
	.A(FE_OFCN47_rank_16_));
   NAND3X1 U819 (.Y(n1515), 
	.C(FE_OFCN165_rank_14_), 
	.B(FE_OFCN166_rank_12_), 
	.A(FE_OFCN167_rank_13_));
   NAND3X1 U820 (.Y(n1519), 
	.C(FE_OFCN176_rank_5_), 
	.B(FE_OFCN177_rank_3_), 
	.A(FE_OFCN178_rank_4_));
   NAND3X1 U821 (.Y(n1526), 
	.C(FE_OFCN2_rank_2_), 
	.B(FE_OFCN0_rank_0_), 
	.A(FE_OFCN1_rank_1_));
   OAI21X1 U822 (.Y(n2050), 
	.C(FE_OFCN308_n1531), 
	.B(n2969), 
	.A(n2831));
   NAND3X1 U823 (.Y(n1531), 
	.C(n2830), 
	.B(n2969), 
	.A(rank[21]));
   OAI21X1 U825 (.Y(n2051), 
	.C(n1535), 
	.B(n1534), 
	.A(rank[21]));
   OAI21X1 U827 (.Y(n2052), 
	.C(FE_OFCN293_n1540), 
	.B(n2872), 
	.A(FE_OFCN294_n1538));
   NAND3X1 U828 (.Y(n1540), 
	.C(n2295), 
	.B(rank[19]), 
	.A(n2842));
   AOI21X1 U830 (.Y(n1538), 
	.C(n1545), 
	.B(n2876), 
	.A(n2842));
   OAI21X1 U831 (.Y(n2053), 
	.C(FE_OFCN292_n1547), 
	.B(n2876), 
	.A(n2843));
   NAND3X1 U832 (.Y(n1547), 
	.C(n2842), 
	.B(n2876), 
	.A(FE_OFCN23_rank_18_));
   OAI21X1 U835 (.Y(n1545), 
	.C(n2379), 
	.B(n1548), 
	.A(FE_OFCN23_rank_18_));
   OAI21X1 U836 (.Y(n2054), 
	.C(n1550), 
	.B(n1548), 
	.A(FE_OFCN23_rank_18_));
   OAI21X1 U838 (.Y(n1548), 
	.C(n2379), 
	.B(n2340), 
	.A(n2946));
   NAND3X1 U841 (.Y(n1553), 
	.C(n1556), 
	.B(n2871), 
	.A(n85));
   NAND3X1 U845 (.Y(n1558), 
	.C(FE_OFCN221_n1561), 
	.B(n2875), 
	.A(n2350));
   AOI21X1 U846 (.Y(n1561), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN24_rank_19_));
   NAND3X1 U848 (.Y(n1557), 
	.C(n88), 
	.B(n2876), 
	.A(n2350));
   OAI21X1 U851 (.Y(n2055), 
	.C(FE_OFCN299_n1567), 
	.B(n2886), 
	.A(FE_OFCN300_n1565));
   NAND3X1 U852 (.Y(n1567), 
	.C(n2294), 
	.B(FE_OFCN47_rank_16_), 
	.A(n2840));
   AOI21X1 U854 (.Y(n1565), 
	.C(n1572), 
	.B(n2888), 
	.A(n2840));
   OAI21X1 U855 (.Y(n2056), 
	.C(FE_OFCN298_n1574), 
	.B(n2888), 
	.A(n2841));
   NAND3X1 U856 (.Y(n1574), 
	.C(n2840), 
	.B(n2888), 
	.A(FE_OFCN46_rank_15_));
   OAI21X1 U859 (.Y(n1572), 
	.C(n2376), 
	.B(n1575), 
	.A(FE_OFCN46_rank_15_));
   OAI21X1 U860 (.Y(n2057), 
	.C(n1577), 
	.B(n1575), 
	.A(FE_OFCN46_rank_15_));
   OAI21X1 U862 (.Y(n1575), 
	.C(n2376), 
	.B(n2336), 
	.A(n2946));
   NAND3X1 U865 (.Y(n1579), 
	.C(n1556), 
	.B(n2968), 
	.A(n84));
   NAND3X1 U869 (.Y(n1582), 
	.C(FE_OFCN219_n1585), 
	.B(n2887), 
	.A(n2349));
   AOI21X1 U870 (.Y(n1585), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN47_rank_16_));
   NAND3X1 U872 (.Y(n1581), 
	.C(n88), 
	.B(n2888), 
	.A(n2349));
   OAI21X1 U875 (.Y(n2058), 
	.C(FE_OFCN296_n1588), 
	.B(n2972), 
	.A(FE_OFCN297_n1586));
   NAND3X1 U876 (.Y(n1588), 
	.C(n2293), 
	.B(rank[13]), 
	.A(n2838));
   AOI21X1 U878 (.Y(n1586), 
	.C(n1593), 
	.B(n2974), 
	.A(n2838));
   OAI21X1 U879 (.Y(n2059), 
	.C(FE_OFCN295_n1595), 
	.B(n2974), 
	.A(n2839));
   NAND3X1 U880 (.Y(n1595), 
	.C(n2838), 
	.B(n2974), 
	.A(rank[12]));
   OAI21X1 U883 (.Y(n1593), 
	.C(n2372), 
	.B(n1596), 
	.A(FE_OFCN166_rank_12_));
   OAI21X1 U884 (.Y(n2060), 
	.C(n1598), 
	.B(n1596), 
	.A(FE_OFCN166_rank_12_));
   OAI21X1 U886 (.Y(n1596), 
	.C(n2372), 
	.B(n2332), 
	.A(n2946));
   NAND3X1 U889 (.Y(n1600), 
	.C(n1556), 
	.B(n2968), 
	.A(n2871));
   NAND3X1 U893 (.Y(n1603), 
	.C(FE_OFCN217_n1606), 
	.B(n2973), 
	.A(n2348));
   AOI21X1 U894 (.Y(n1606), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN167_rank_13_));
   NAND3X1 U896 (.Y(n1602), 
	.C(n88), 
	.B(n2974), 
	.A(n2348));
   OAI21X1 U899 (.Y(n2061), 
	.C(FE_OFCN311_n1609), 
	.B(n2978), 
	.A(FE_OFCN312_n1607));
   NAND3X1 U900 (.Y(n1609), 
	.C(n2292), 
	.B(FE_OFCN174_rank_10_), 
	.A(n2836));
   AOI21X1 U902 (.Y(n1607), 
	.C(n1614), 
	.B(n2980), 
	.A(n2836));
   OAI21X1 U903 (.Y(n2062), 
	.C(FE_OFCN310_n1616), 
	.B(n2980), 
	.A(n2837));
   NAND3X1 U904 (.Y(n1616), 
	.C(n2836), 
	.B(n2980), 
	.A(rank[9]));
   OAI21X1 U907 (.Y(n1614), 
	.C(n2369), 
	.B(n1617), 
	.A(rank[9]));
   OAI21X1 U908 (.Y(n2063), 
	.C(n1619), 
	.B(n1617), 
	.A(FE_OFCN173_rank_9_));
   OAI21X1 U910 (.Y(n1617), 
	.C(n2369), 
	.B(n2328), 
	.A(n2946));
   NAND3X1 U913 (.Y(n1621), 
	.C(n1623), 
	.B(n84), 
	.A(n85));
   NAND3X1 U917 (.Y(n1625), 
	.C(FE_OFCN215_n1628), 
	.B(n2979), 
	.A(n2347));
   AOI21X1 U918 (.Y(n1628), 
	.C(n89), 
	.B(n2773), 
	.A(rank[10]));
   NAND3X1 U920 (.Y(n1624), 
	.C(n88), 
	.B(n2980), 
	.A(n2347));
   OAI21X1 U923 (.Y(n2064), 
	.C(FE_OFCN305_n1631), 
	.B(n2975), 
	.A(FE_OFCN306_n1629));
   NAND3X1 U924 (.Y(n1631), 
	.C(n2291), 
	.B(rank[7]), 
	.A(n2834));
   AOI21X1 U926 (.Y(n1629), 
	.C(n1636), 
	.B(n2977), 
	.A(n2834));
   OAI21X1 U927 (.Y(n2065), 
	.C(FE_OFCN304_n1638), 
	.B(n2977), 
	.A(n2835));
   NAND3X1 U928 (.Y(n1638), 
	.C(n2834), 
	.B(n2977), 
	.A(rank[6]));
   OAI21X1 U931 (.Y(n1636), 
	.C(n2366), 
	.B(n1639), 
	.A(rank[6]));
   OAI21X1 U932 (.Y(n2066), 
	.C(n1641), 
	.B(n1639), 
	.A(FE_OFCN170_rank_6_));
   OAI21X1 U934 (.Y(n1639), 
	.C(n2366), 
	.B(n2324), 
	.A(n2946));
   NAND3X1 U937 (.Y(n1643), 
	.C(n1623), 
	.B(n2871), 
	.A(n85));
   NAND3X1 U941 (.Y(n1646), 
	.C(FE_OFCN213_n1649), 
	.B(n2976), 
	.A(n2564));
   AOI21X1 U942 (.Y(n1649), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN171_rank_7_));
   NAND3X1 U944 (.Y(n1645), 
	.C(n88), 
	.B(n2977), 
	.A(n2564));
   OAI21X1 U947 (.Y(n2067), 
	.C(FE_OFCN302_n1652), 
	.B(n2981), 
	.A(FE_OFCN303_n1650));
   NAND3X1 U948 (.Y(n1652), 
	.C(n2290), 
	.B(rank[4]), 
	.A(n2832));
   AOI21X1 U950 (.Y(n1650), 
	.C(n1657), 
	.B(n2983), 
	.A(n2832));
   OAI21X1 U951 (.Y(n2068), 
	.C(FE_OFCN301_n1659), 
	.B(n2983), 
	.A(n2833));
   NAND3X1 U952 (.Y(n1659), 
	.C(n2832), 
	.B(n2983), 
	.A(FE_OFCN177_rank_3_));
   OAI21X1 U955 (.Y(n1657), 
	.C(n2362), 
	.B(n1660), 
	.A(FE_OFCN177_rank_3_));
   OAI21X1 U956 (.Y(n2069), 
	.C(n1662), 
	.B(n1660), 
	.A(FE_OFCN177_rank_3_));
   OAI21X1 U958 (.Y(n1660), 
	.C(n2362), 
	.B(n2320), 
	.A(n2946));
   NAND3X1 U961 (.Y(n1664), 
	.C(n1623), 
	.B(n2968), 
	.A(n84));
   NAND3X1 U965 (.Y(n1667), 
	.C(FE_OFCN224_n1670), 
	.B(n2982), 
	.A(n2346));
   AOI21X1 U966 (.Y(n1670), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN178_rank_4_));
   NAND3X1 U968 (.Y(n1666), 
	.C(n88), 
	.B(n2983), 
	.A(n2346));
   OAI21X1 U971 (.Y(n2070), 
	.C(FE_OFCN314_n1673), 
	.B(n2850), 
	.A(FE_OFCN315_n1671));
   NAND3X1 U972 (.Y(n1673), 
	.C(n2289), 
	.B(FE_OFCN1_rank_1_), 
	.A(n2828));
   AOI21X1 U974 (.Y(n1671), 
	.C(n1678), 
	.B(n2849), 
	.A(n2828));
   OAI21X1 U975 (.Y(n2071), 
	.C(FE_OFCN313_n1680), 
	.B(n2849), 
	.A(n2829));
   NAND3X1 U976 (.Y(n1680), 
	.C(n2828), 
	.B(n2849), 
	.A(FE_OFCN0_rank_0_));
   OAI21X1 U979 (.Y(n1678), 
	.C(n2354), 
	.B(n1681), 
	.A(FE_OFCN0_rank_0_));
   OAI21X1 U980 (.Y(n2072), 
	.C(FE_OFCN307_n1685), 
	.B(n2971), 
	.A(FE_OFCN309_n1683));
   NAND3X1 U981 (.Y(n1685), 
	.C(n2288), 
	.B(rank[22]), 
	.A(n2830));
   AOI21X1 U983 (.Y(n1683), 
	.C(n1533), 
	.B(n2969), 
	.A(n2830));
   OAI21X1 U984 (.Y(n1533), 
	.C(n2358), 
	.B(n1534), 
	.A(FE_OFCN163_rank_21_));
   OAI21X1 U986 (.Y(n1534), 
	.C(n2358), 
	.B(n2316), 
	.A(n2946));
   NAND3X1 U989 (.Y(n1688), 
	.C(n1556), 
	.B(n84), 
	.A(n85));
   NOR3X1 U990 (.Y(n1556), 
	.C(n2885), 
	.B(j_3_), 
	.A(n2752));
   NAND3X1 U995 (.Y(n1691), 
	.C(FE_OFCN211_n1694), 
	.B(n2970), 
	.A(n2345));
   AOI21X1 U996 (.Y(n1694), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN162_rank_22_));
   NAND3X1 U998 (.Y(n1690), 
	.C(n88), 
	.B(n2969), 
	.A(n2345));
   OAI21X1 U1001 (.Y(n2073), 
	.C(n1695), 
	.B(n1681), 
	.A(rank[0]));
   OAI21X1 U1003 (.Y(n1681), 
	.C(n2354), 
	.B(n2312), 
	.A(n2946));
   NAND3X1 U1010 (.Y(n1697), 
	.C(n1623), 
	.B(n2968), 
	.A(n2871));
   NOR3X1 U1011 (.Y(n1623), 
	.C(n2752), 
	.B(n86), 
	.A(j_3_));
   NAND3X1 U1018 (.Y(n1700), 
	.C(FE_OFCN209_n1703), 
	.B(n2845), 
	.A(n2344));
   AOI21X1 U1019 (.Y(n1703), 
	.C(n89), 
	.B(n2773), 
	.A(FE_OFCN1_rank_1_));
   NAND3X1 U1023 (.Y(n1699), 
	.C(n88), 
	.B(n2849), 
	.A(n2344));
   AND2X1 U1209 (.Y(n1212), 
	.B(DIN[12]), 
	.A(mem[20]));
   AND2X1 U1210 (.Y(n1163), 
	.B(DIN[9]), 
	.A(FE_OFCN122_mem_81_));
   AND2X1 U1211 (.Y(n1099), 
	.B(DIN[9]), 
	.A(FE_OFCN42_mem_113_));
   AND2X1 U1212 (.Y(n1083), 
	.B(DIN[11]), 
	.A(FE_OFCN40_mem_115_));
   AND2X1 U1213 (.Y(n1292), 
	.B(DIN[9]), 
	.A(mem[49]));
   AND2X1 U1214 (.Y(n1524), 
	.B(FE_OFCN199_n1520), 
	.A(FE_OFCN198_n1521));
   AND2X1 U1215 (.Y(n905), 
	.B(n2537), 
	.A(FE_OFCN250_n1005));
   OR2X1 U1216 (.Y(n1662), 
	.B(n2982), 
	.A(n2362));
   OR2X1 U1217 (.Y(n1619), 
	.B(n2979), 
	.A(n2369));
   OR2X1 U1218 (.Y(n1641), 
	.B(n2976), 
	.A(n2366));
   OR2X1 U1219 (.Y(n1598), 
	.B(n2973), 
	.A(n2372));
   OR2X1 U1220 (.Y(n1535), 
	.B(n2970), 
	.A(n2358));
   AND2X1 U1221 (.Y(n1781), 
	.B(n2557), 
	.A(n2752));
   AND2X1 U1222 (.Y(n874), 
	.B(n2827), 
	.A(match));
   OR2X1 U1223 (.Y(n1577), 
	.B(n2887), 
	.A(n2376));
   OR2X1 U1224 (.Y(n1550), 
	.B(n2875), 
	.A(n2379));
   OR2X1 U1225 (.Y(n1695), 
	.B(n2845), 
	.A(n2354));
   OR2X1 U1226 (.Y(n904), 
	.B(n2730), 
	.A(n2844));
   AND2X1 U1227 (.Y(n868), 
	.B(EN), 
	.A(m));
   AND2X1 U1228 (.Y(n1003), 
	.B(n1018), 
	.A(n1017));
   AND2X1 U1229 (.Y(n1528), 
	.B(FE_OFCN195_n1513), 
	.A(FE_OFCN183_n1522));
   OR2X1 U1230 (.Y(n878), 
	.B(WE), 
	.A(n2666));
   OR2X1 U1292 (.Y(n2312), 
	.B(n2315), 
	.A(n2314));
   OR2X1 U1293 (.Y(n2315), 
	.B(n2313), 
	.A(n1701));
   OR2X1 U1294 (.Y(n2316), 
	.B(n2319), 
	.A(n2318));
   OR2X1 U1295 (.Y(n2319), 
	.B(n2317), 
	.A(n1692));
   OR2X1 U1296 (.Y(n2320), 
	.B(n2323), 
	.A(n2322));
   OR2X1 U1297 (.Y(n2323), 
	.B(n2321), 
	.A(n1668));
   OR2X1 U1298 (.Y(n2324), 
	.B(n2327), 
	.A(n2326));
   OR2X1 U1299 (.Y(n2327), 
	.B(n2325), 
	.A(n1647));
   OR2X1 U1300 (.Y(n2328), 
	.B(n2331), 
	.A(n2330));
   OR2X1 U1301 (.Y(n2331), 
	.B(n2329), 
	.A(n1626));
   OR2X1 U1302 (.Y(n2332), 
	.B(n2335), 
	.A(n2334));
   OR2X1 U1303 (.Y(n2335), 
	.B(n2333), 
	.A(n1604));
   OR2X1 U1304 (.Y(n2336), 
	.B(n2339), 
	.A(n2338));
   OR2X1 U1305 (.Y(n2339), 
	.B(n2337), 
	.A(n1583));
   OR2X1 U1306 (.Y(n2340), 
	.B(n2343), 
	.A(n2342));
   OR2X1 U1307 (.Y(n2343), 
	.B(n2341), 
	.A(n1559));
   OR2X1 U1308 (.Y(n2354), 
	.B(n2357), 
	.A(n2356));
   OR2X1 U1309 (.Y(n2357), 
	.B(n2355), 
	.A(n1698));
   OR2X1 U1310 (.Y(n2358), 
	.B(n2361), 
	.A(n2360));
   OR2X1 U1311 (.Y(n2361), 
	.B(n2359), 
	.A(n1689));
   OR2X1 U1312 (.Y(n2362), 
	.B(n2365), 
	.A(n2364));
   OR2X1 U1313 (.Y(n2365), 
	.B(n2363), 
	.A(n1665));
   OR2X1 U1314 (.Y(n2366), 
	.B(n2368), 
	.A(n2367));
   OR2X1 U1315 (.Y(n2368), 
	.B(n2359), 
	.A(n1644));
   OR2X1 U1316 (.Y(n2369), 
	.B(n2371), 
	.A(n2370));
   OR2X1 U1317 (.Y(n2371), 
	.B(n2355), 
	.A(n1622));
   OR2X1 U1318 (.Y(n2372), 
	.B(n2375), 
	.A(n2374));
   OR2X1 U1319 (.Y(n2375), 
	.B(n2373), 
	.A(n1601));
   OR2X1 U1320 (.Y(n2376), 
	.B(n2378), 
	.A(n2377));
   OR2X1 U1321 (.Y(n2378), 
	.B(n2363), 
	.A(n1580));
   OR2X1 U1322 (.Y(n2379), 
	.B(n2381), 
	.A(n2380));
   OR2X1 U1323 (.Y(n2381), 
	.B(n2373), 
	.A(n1554));
   AND2X1 U1324 (.Y(n2989), 
	.B(n2815), 
	.A(n2818));
   AND2X1 U1325 (.Y(n1701), 
	.B(n2850), 
	.A(n87));
   AND2X1 U1326 (.Y(n1698), 
	.B(n2312), 
	.A(n868));
   AND2X1 U1327 (.Y(n1692), 
	.B(n2971), 
	.A(n87));
   AND2X1 U1328 (.Y(n1689), 
	.B(n2316), 
	.A(n868));
   AND2X1 U1329 (.Y(n1668), 
	.B(n2981), 
	.A(n87));
   AND2X1 U1330 (.Y(n1665), 
	.B(n2320), 
	.A(n868));
   AND2X1 U1331 (.Y(n1647), 
	.B(n2975), 
	.A(n87));
   AND2X1 U1332 (.Y(n1644), 
	.B(n2324), 
	.A(n868));
   AND2X1 U1333 (.Y(n1626), 
	.B(n2978), 
	.A(n87));
   AND2X1 U1334 (.Y(n1622), 
	.B(n2328), 
	.A(n868));
   AND2X1 U1335 (.Y(n1604), 
	.B(n2972), 
	.A(n87));
   AND2X1 U1336 (.Y(n1601), 
	.B(n2332), 
	.A(n868));
   AND2X1 U1337 (.Y(n1583), 
	.B(n2886), 
	.A(n87));
   AND2X1 U1338 (.Y(n1580), 
	.B(n2336), 
	.A(n868));
   AND2X1 U1339 (.Y(n1559), 
	.B(n2872), 
	.A(n87));
   AND2X1 U1340 (.Y(n1554), 
	.B(n2340), 
	.A(n868));
   AND2X1 U1372 (.Y(n1504), 
	.B(DIN[5]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1373 (.Y(n2166), 
	.A(n1504));
   AND2X1 U1374 (.Y(n1499), 
	.B(n1314), 
	.A(FE_OFCN288_n1485));
   INVX1 U1375 (.Y(n2167), 
	.A(n1499));
   AND2X1 U1376 (.Y(n1498), 
	.B(n1312), 
	.A(FE_OFCN288_n1485));
   INVX1 U1377 (.Y(n2168), 
	.A(n1498));
   AND2X1 U1378 (.Y(n1497), 
	.B(n1310), 
	.A(FE_OFCN288_n1485));
   INVX1 U1379 (.Y(n2169), 
	.A(n1497));
   AND2X1 U1380 (.Y(n1496), 
	.B(n1308), 
	.A(FE_OFCN288_n1485));
   INVX1 U1381 (.Y(n2170), 
	.A(n1496));
   AND2X1 U1382 (.Y(n1488), 
	.B(n250), 
	.A(FE_OFCN288_n1485));
   INVX1 U1383 (.Y(n2171), 
	.A(n1488));
   AND2X1 U1384 (.Y(n1487), 
	.B(n251), 
	.A(FE_OFCN288_n1485));
   INVX1 U1385 (.Y(n2172), 
	.A(n1487));
   AND2X1 U1386 (.Y(n1486), 
	.B(n252), 
	.A(FE_OFCN288_n1485));
   INVX1 U1387 (.Y(n2173), 
	.A(n1486));
   AND2X1 U1388 (.Y(n1475), 
	.B(FE_OFCN317_n1463), 
	.A(mem[23]));
   INVX1 U1389 (.Y(n2174), 
	.A(n1475));
   AND2X1 U1390 (.Y(n1473), 
	.B(FE_OFCN317_n1463), 
	.A(mem[25]));
   INVX1 U1391 (.Y(n2175), 
	.A(n1473));
   AND2X1 U1392 (.Y(n1472), 
	.B(FE_OFCN317_n1463), 
	.A(mem[26]));
   INVX1 U1393 (.Y(n2176), 
	.A(n1472));
   AND2X1 U1394 (.Y(n1471), 
	.B(FE_OFCN317_n1463), 
	.A(mem[27]));
   INVX1 U1395 (.Y(n2177), 
	.A(n1471));
   AND2X1 U1396 (.Y(n1470), 
	.B(FE_OFCN317_n1463), 
	.A(mem[28]));
   INVX1 U1397 (.Y(n2178), 
	.A(n1470));
   AND2X1 U1398 (.Y(n1467), 
	.B(FE_OFCN317_n1463), 
	.A(mem[31]));
   INVX1 U1399 (.Y(n2179), 
	.A(n1467));
   AND2X1 U1400 (.Y(n1466), 
	.B(n1463), 
	.A(matchN[3]));
   INVX1 U1401 (.Y(n2180), 
	.A(n1466));
   AND2X2 U1402 (.Y(n1465), 
	.B(n1463), 
	.A(matchN[4]));
   INVX1 U1403 (.Y(n2181), 
	.A(n1465));
   AND2X1 U1404 (.Y(n1464), 
	.B(n1463), 
	.A(matchN[5]));
   INVX1 U1405 (.Y(n2182), 
	.A(n1464));
   AND2X1 U1406 (.Y(n1462), 
	.B(DIN[0]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1407 (.Y(n2183), 
	.A(n1462));
   AND2X1 U1408 (.Y(n1461), 
	.B(DIN[1]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1409 (.Y(n2184), 
	.A(n1461));
   AND2X1 U1410 (.Y(n1460), 
	.B(DIN[2]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1411 (.Y(n2185), 
	.A(n1460));
   AND2X1 U1412 (.Y(n1459), 
	.B(DIN[3]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1413 (.Y(n2186), 
	.A(n1459));
   AND2X1 U1414 (.Y(n1458), 
	.B(DIN[4]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1415 (.Y(n2187), 
	.A(n1458));
   AND2X1 U1416 (.Y(n1453), 
	.B(DIN[7]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1417 (.Y(n2188), 
	.A(n1453));
   AND2X1 U1418 (.Y(n1452), 
	.B(n1314), 
	.A(n1437));
   INVX1 U1419 (.Y(n2189), 
	.A(n1452));
   AND2X1 U1420 (.Y(n1433), 
	.B(FE_OFCN318_n1417), 
	.A(mem[51]));
   INVX1 U1421 (.Y(n2190), 
	.A(n1433));
   AND2X1 U1422 (.Y(n1432), 
	.B(FE_OFCN318_n1417), 
	.A(FE_OFCN138_mem_52_));
   INVX1 U1423 (.Y(n2191), 
	.A(n1432));
   AND2X1 U1424 (.Y(n1426), 
	.B(FE_OFCN318_n1417), 
	.A(FE_OFCN132_mem_58_));
   INVX1 U1425 (.Y(n2192), 
	.A(n1426));
   AND2X1 U1426 (.Y(n1425), 
	.B(FE_OFCN318_n1417), 
	.A(mem[59]));
   INVX1 U1427 (.Y(n2193), 
	.A(n1425));
   AND2X1 U1428 (.Y(n1424), 
	.B(FE_OFCN318_n1417), 
	.A(mem[60]));
   INVX1 U1429 (.Y(n2194), 
	.A(n1424));
   AND2X1 U1430 (.Y(n1422), 
	.B(FE_OFCN318_n1417), 
	.A(FE_OFCN128_mem_62_));
   INVX1 U1431 (.Y(n2195), 
	.A(n1422));
   AND2X1 U1432 (.Y(n1421), 
	.B(FE_OFCN318_n1417), 
	.A(mem[63]));
   INVX1 U1433 (.Y(n2196), 
	.A(n1421));
   AND2X1 U1434 (.Y(n1420), 
	.B(n1417), 
	.A(matchN[9]));
   INVX1 U1435 (.Y(n2197), 
	.A(n1420));
   AND2X1 U1436 (.Y(n1419), 
	.B(n1417), 
	.A(FE_OFCN125_matchN_10_));
   INVX1 U1437 (.Y(n2198), 
	.A(n1419));
   AND2X1 U1438 (.Y(n1418), 
	.B(n1417), 
	.A(matchN[11]));
   INVX1 U1439 (.Y(n2199), 
	.A(n1418));
   AND2X1 U1440 (.Y(n1416), 
	.B(DIN[0]), 
	.A(n1391));
   INVX1 U1441 (.Y(n2200), 
	.A(n1416));
   AND2X1 U1442 (.Y(n1415), 
	.B(DIN[1]), 
	.A(n1391));
   INVX1 U1443 (.Y(n2201), 
	.A(n1415));
   AND2X1 U1444 (.Y(n1414), 
	.B(DIN[2]), 
	.A(n1391));
   INVX1 U1445 (.Y(n2202), 
	.A(n1414));
   AND2X1 U1446 (.Y(n1413), 
	.B(DIN[3]), 
	.A(FE_OFCN290_n1391));
   INVX1 U1447 (.Y(n2203), 
	.A(n1413));
   AND2X1 U1448 (.Y(n1407), 
	.B(DIN[7]), 
	.A(FE_OFCN290_n1391));
   INVX1 U1449 (.Y(n2204), 
	.A(n1407));
   AND2X1 U1450 (.Y(n1406), 
	.B(n1314), 
	.A(n1391));
   INVX1 U1451 (.Y(n2205), 
	.A(n1406));
   AND2X1 U1452 (.Y(n1405), 
	.B(n1312), 
	.A(FE_OFCN290_n1391));
   INVX1 U1453 (.Y(n2206), 
	.A(n1405));
   AND2X1 U1454 (.Y(n1404), 
	.B(n1310), 
	.A(n1391));
   INVX1 U1455 (.Y(n2207), 
	.A(n1404));
   AND2X1 U1456 (.Y(n1387), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN120_mem_83_));
   INVX1 U1457 (.Y(n2208), 
	.A(n1387));
   AND2X1 U1458 (.Y(n1386), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN119_mem_84_));
   INVX1 U1459 (.Y(n2209), 
	.A(n1386));
   AND2X1 U1460 (.Y(n1382), 
	.B(n1371), 
	.A(mem[88]));
   INVX1 U1461 (.Y(n2210), 
	.A(n1382));
   AND2X1 U1462 (.Y(n1379), 
	.B(FE_OFCN319_n1371), 
	.A(mem[91]));
   INVX1 U1463 (.Y(n2211), 
	.A(n1379));
   AND2X1 U1464 (.Y(n1378), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN111_mem_92_));
   INVX1 U1465 (.Y(n2212), 
	.A(n1378));
   AND2X1 U1466 (.Y(n1376), 
	.B(FE_OFCN319_n1371), 
	.A(mem[94]));
   INVX1 U1467 (.Y(n2213), 
	.A(n1376));
   AND2X1 U1468 (.Y(n1375), 
	.B(FE_OFCN319_n1371), 
	.A(mem[95]));
   INVX1 U1469 (.Y(n2214), 
	.A(n1375));
   AND2X1 U1470 (.Y(n1374), 
	.B(n1371), 
	.A(FE_OFCN107_matchN_15_));
   INVX1 U1471 (.Y(n2215), 
	.A(n1374));
   AND2X1 U1472 (.Y(n1373), 
	.B(n1371), 
	.A(FE_OFCN106_matchN_16_));
   INVX1 U1473 (.Y(n2216), 
	.A(n1373));
   AND2X1 U1474 (.Y(n1372), 
	.B(n1371), 
	.A(matchN[17]));
   INVX1 U1475 (.Y(n2217), 
	.A(n1372));
   AND2X1 U1476 (.Y(n1356), 
	.B(n1314), 
	.A(FE_OFCN291_n1335));
   INVX1 U1477 (.Y(n2218), 
	.A(n1356));
   AND2X1 U1478 (.Y(n1354), 
	.B(n1312), 
	.A(FE_OFCN291_n1335));
   INVX1 U1479 (.Y(n2219), 
	.A(n1354));
   AND2X1 U1480 (.Y(n1352), 
	.B(n1310), 
	.A(FE_OFCN291_n1335));
   INVX1 U1481 (.Y(n2220), 
	.A(n1352));
   AND2X1 U1482 (.Y(n1350), 
	.B(n1308), 
	.A(FE_OFCN291_n1335));
   INVX1 U1483 (.Y(n2221), 
	.A(n1350));
   AND2X1 U1484 (.Y(n1339), 
	.B(n1300), 
	.A(FE_OFCN291_n1335));
   INVX1 U1485 (.Y(n2222), 
	.A(n1339));
   AND2X1 U1486 (.Y(n1337), 
	.B(n251), 
	.A(FE_OFCN291_n1335));
   INVX1 U1487 (.Y(n2223), 
	.A(n1337));
   AND2X1 U1488 (.Y(n1336), 
	.B(n252), 
	.A(FE_OFCN291_n1335));
   INVX1 U1489 (.Y(n2224), 
	.A(n1336));
   AND2X1 U1490 (.Y(n1325), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN40_mem_115_));
   INVX1 U1491 (.Y(n2225), 
	.A(n1325));
   AND2X1 U1492 (.Y(n1323), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN39_mem_116_));
   INVX1 U1493 (.Y(n2226), 
	.A(n1323));
   AND2X1 U1494 (.Y(n1315), 
	.B(FE_OFCN320_n1021), 
	.A(mem[120]));
   INVX1 U1495 (.Y(n2227), 
	.A(n1315));
   AND2X1 U1496 (.Y(n1313), 
	.B(FE_OFCN320_n1021), 
	.A(mem[121]));
   INVX1 U1497 (.Y(n2228), 
	.A(n1313));
   AND2X1 U1498 (.Y(n1309), 
	.B(FE_OFCN320_n1021), 
	.A(mem[123]));
   INVX1 U1499 (.Y(n2229), 
	.A(n1309));
   AND2X1 U1500 (.Y(n1307), 
	.B(FE_OFCN320_n1021), 
	.A(mem[124]));
   INVX1 U1501 (.Y(n2230), 
	.A(n1307));
   AND2X1 U1502 (.Y(n1303), 
	.B(FE_OFCN320_n1021), 
	.A(mem[126]));
   INVX1 U1503 (.Y(n2231), 
	.A(n1303));
   AND2X1 U1504 (.Y(n1301), 
	.B(FE_OFCN320_n1021), 
	.A(mem[127]));
   INVX1 U1505 (.Y(n2232), 
	.A(n1301));
   AND2X1 U1506 (.Y(n1036), 
	.B(n1037), 
	.A(n1028));
   INVX1 U1507 (.Y(n2233), 
	.A(n1036));
   AND2X1 U1508 (.Y(n1033), 
	.B(FE_OFCN201_n1034), 
	.A(n1028));
   INVX1 U1509 (.Y(n2234), 
	.A(n1033));
   AND2X1 U1510 (.Y(n1030), 
	.B(FE_OFCN197_n1031), 
	.A(n1028));
   INVX1 U1511 (.Y(n2235), 
	.A(n1030));
   AND2X1 U1512 (.Y(n1025), 
	.B(n1021), 
	.A(FE_OFCN26_matchN_22_));
   INVX1 U1513 (.Y(n2236), 
	.A(n1025));
   AND2X1 U1514 (.Y(n1023), 
	.B(n1021), 
	.A(FE_OFCN25_matchN_23_));
   INVX1 U1515 (.Y(n2237), 
	.A(n1023));
   AND2X1 U1516 (.Y(n990), 
	.B(FE_PSN325_n991), 
	.A(n897));
   INVX2 U1517 (.Y(n2238), 
	.A(n990));
   AND2X1 U1518 (.Y(n987), 
	.B(n897), 
	.A(FE_OFCN251_n988));
   INVX2 U1519 (.Y(n2239), 
	.A(n987));
   AND2X1 U1520 (.Y(n974), 
	.B(FE_PSN323_n975), 
	.A(n906));
   INVX2 U1521 (.Y(n2240), 
	.A(n974));
   AND2X1 U1522 (.Y(n959), 
	.B(FE_PSN330_n960), 
	.A(FE_OFCN261_n888));
   INVX2 U1523 (.Y(n2241), 
	.A(n959));
   AND2X1 U1524 (.Y(n956), 
	.B(FE_PSN332_FE_OFCN261_n888), 
	.A(n957));
   INVX2 U1525 (.Y(n2242), 
	.A(n956));
   AND2X1 U1526 (.Y(n943), 
	.B(n944), 
	.A(FE_OFCN263_n886));
   INVX2 U1527 (.Y(n2243), 
	.A(n943));
   AND2X1 U1528 (.Y(n925), 
	.B(FE_PSN324_n926), 
	.A(FE_OFCN268_n892));
   INVX2 U1529 (.Y(n2244), 
	.A(n925));
   OR2X2 U1531 (.Y(n971), 
	.B(n2808), 
	.A(n972));
   INVX2 U1532 (.Y(n2246), 
	.A(n971));
   OR2X2 U1533 (.Y(n940), 
	.B(n2804), 
	.A(n941));
   INVX2 U1534 (.Y(n2247), 
	.A(n940));
   AND2X1 U1537 (.Y(n986), 
	.B(n975), 
	.A(n2955));
   INVX1 U1538 (.Y(n2250), 
	.A(n986));
   AND2X2 U1539 (.Y(n955), 
	.B(n944), 
	.A(n2948));
   INVX2 U1540 (.Y(n2251), 
	.A(n955));
   AND2X1 U1541 (.Y(n915), 
	.B(FE_OFCN27_matchN_21_), 
	.A(n2799));
   INVX2 U1542 (.Y(n2252), 
	.A(n915));
   AND2X1 U1557 (.Y(n1016), 
	.B(n2854), 
	.A(matchN[3]));
   INVX2 U1558 (.Y(n2267), 
	.A(n1016));
   AND2X1 U1559 (.Y(n1001), 
	.B(n991), 
	.A(n2926));
   INVX4 U1560 (.Y(n2268), 
	.A(n1001));
   AND2X2 U1561 (.Y(n970), 
	.B(n960), 
	.A(n2907));
   INVX2 U1562 (.Y(n2269), 
	.A(n970));
   AND2X2 U1563 (.Y(n939), 
	.B(n926), 
	.A(n2929));
   INVX2 U1564 (.Y(n2270), 
	.A(n939));
   OR2X1 U1582 (.Y(n1686), 
	.B(n2970), 
	.A(FE_OFCN164_rank_23_));
   INVX1 U1583 (.Y(n2288), 
	.A(n1686));
   OR2X1 U1584 (.Y(n1675), 
	.B(n2845), 
	.A(FE_OFCN2_rank_2_));
   INVX1 U1585 (.Y(n2289), 
	.A(n1675));
   OR2X1 U1586 (.Y(n1654), 
	.B(n2982), 
	.A(rank[5]));
   INVX1 U1587 (.Y(n2290), 
	.A(n1654));
   OR2X1 U1588 (.Y(n1633), 
	.B(n2976), 
	.A(rank[8]));
   INVX1 U1589 (.Y(n2291), 
	.A(n1633));
   OR2X1 U1590 (.Y(n1611), 
	.B(n2979), 
	.A(rank[11]));
   INVX1 U1591 (.Y(n2292), 
	.A(n1611));
   OR2X1 U1592 (.Y(n1590), 
	.B(n2973), 
	.A(rank[14]));
   INVX1 U1593 (.Y(n2293), 
	.A(n1590));
   OR2X1 U1594 (.Y(n1569), 
	.B(n2887), 
	.A(rank[17]));
   INVX1 U1595 (.Y(n2294), 
	.A(n1569));
   OR2X1 U1596 (.Y(n1542), 
	.B(n2875), 
	.A(rank[20]));
   INVX1 U1597 (.Y(n2295), 
	.A(n1542));
   OR2X1 U1598 (.Y(n1527), 
	.B(n2351), 
	.A(FE_OFCN197_n1031));
   INVX1 U1599 (.Y(n2296), 
	.A(n1527));
   OR2X1 U1600 (.Y(n1257), 
	.B(mem[37]), 
	.A(mem[38]));
   INVX1 U1601 (.Y(n2297), 
	.A(n1257));
   OR2X2 U1602 (.Y(n1193), 
	.B(mem[6]), 
	.A(mem[7]));
   INVX2 U1603 (.Y(n2298), 
	.A(n1193));
   OR2X1 U1604 (.Y(n1171), 
	.B(n1017), 
	.A(n1011));
   INVX1 U1605 (.Y(n2299), 
	.A(n1171));
   OR2X1 U1606 (.Y(n1128), 
	.B(mem[69]), 
	.A(FE_OFCN54_mem_70_));
   INVX1 U1607 (.Y(n2300), 
	.A(n1128));
   OR2X1 U1608 (.Y(n1064), 
	.B(FE_OFCN97_mem_101_), 
	.A(FE_OFCN96_mem_102_));
   INVX1 U1609 (.Y(n2301), 
	.A(n1064));
   BUFX2 U1611 (.Y(match), 
	.A(FE_OFCN104_n2999));
   INVX1 U1612 (.Y(n2304), 
	.A(FE_OFCN198_n1521));
   INVX1 U1617 (.Y(n2309), 
	.A(matchN[18]));
   INVX1 U1620 (.Y(n2313), 
	.A(FE_OFCN210_n1700));
   INVX1 U1621 (.Y(n2314), 
	.A(FE_OFCN202_n1699));
   INVX1 U1622 (.Y(n2317), 
	.A(FE_OFCN212_n1691));
   INVX1 U1623 (.Y(n2318), 
	.A(FE_OFCN203_n1690));
   INVX1 U1624 (.Y(n2321), 
	.A(FE_OFCN225_n1667));
   INVX1 U1625 (.Y(n2322), 
	.A(FE_OFCN223_n1666));
   INVX1 U1626 (.Y(n2325), 
	.A(FE_OFCN214_n1646));
   INVX1 U1627 (.Y(n2326), 
	.A(FE_OFCN204_n1645));
   INVX1 U1628 (.Y(n2329), 
	.A(FE_OFCN216_n1625));
   INVX1 U1629 (.Y(n2330), 
	.A(FE_OFCN205_n1624));
   INVX1 U1630 (.Y(n2333), 
	.A(FE_OFCN218_n1603));
   INVX1 U1631 (.Y(n2334), 
	.A(FE_OFCN206_n1602));
   INVX1 U1632 (.Y(n2337), 
	.A(FE_OFCN220_n1582));
   INVX1 U1633 (.Y(n2338), 
	.A(FE_OFCN207_n1581));
   INVX1 U1634 (.Y(n2341), 
	.A(FE_OFCN222_n1558));
   INVX1 U1635 (.Y(n2342), 
	.A(FE_OFCN208_n1557));
   AND2X1 U1636 (.Y(n1702), 
	.B(n2774), 
	.A(FE_OFCN2_rank_2_));
   INVX1 U1637 (.Y(n2344), 
	.A(n1702));
   AND2X1 U1638 (.Y(n1693), 
	.B(n2774), 
	.A(FE_OFCN164_rank_23_));
   INVX1 U1639 (.Y(n2345), 
	.A(n1693));
   AND2X1 U1640 (.Y(n1669), 
	.B(n2774), 
	.A(rank[5]));
   INVX1 U1641 (.Y(n2346), 
	.A(n1669));
   AND2X1 U1642 (.Y(n1627), 
	.B(n2774), 
	.A(rank[11]));
   INVX1 U1643 (.Y(n2347), 
	.A(n1627));
   AND2X1 U1644 (.Y(n1605), 
	.B(n2774), 
	.A(rank[14]));
   INVX1 U1645 (.Y(n2348), 
	.A(n1605));
   AND2X1 U1646 (.Y(n1584), 
	.B(n2774), 
	.A(rank[17]));
   INVX1 U1647 (.Y(n2349), 
	.A(n1584));
   AND2X1 U1648 (.Y(n1560), 
	.B(n2774), 
	.A(FE_OFCN22_rank_20_));
   INVX1 U1649 (.Y(n2350), 
	.A(n1560));
   INVX1 U1650 (.Y(n2351), 
	.A(n1524));
   INVX1 U1653 (.Y(n2355), 
	.A(n904));
   INVX1 U1654 (.Y(n2356), 
	.A(FE_OFCN280_n1697));
   INVX1 U1655 (.Y(n2359), 
	.A(n904));
   INVX1 U1656 (.Y(n2360), 
	.A(FE_OFCN284_n1688));
   INVX1 U1657 (.Y(n2363), 
	.A(n904));
   INVX1 U1658 (.Y(n2364), 
	.A(FE_OFCN281_n1664));
   INVX1 U1659 (.Y(n2367), 
	.A(FE_OFCN282_n1643));
   INVX1 U1660 (.Y(n2370), 
	.A(FE_OFCN283_n1621));
   INVX1 U1661 (.Y(n2373), 
	.A(n904));
   INVX1 U1662 (.Y(n2374), 
	.A(FE_OFCN285_n1600));
   INVX1 U1663 (.Y(n2377), 
	.A(FE_OFCN286_n1579));
   INVX1 U1664 (.Y(n2380), 
	.A(FE_OFCN287_n1553));
   INVX1 U1666 (.Y(n2383), 
	.A(FE_OFCN185_n1517));
   AND2X1 U1669 (.Y(n1505), 
	.B(DIN[4]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1670 (.Y(n2386), 
	.A(n1505));
   AND2X1 U1671 (.Y(n1311), 
	.B(FE_OFCN320_n1021), 
	.A(mem[122]));
   INVX1 U1672 (.Y(n2387), 
	.A(n1311));
   AND2X1 U1673 (.Y(n879), 
	.B(n2666), 
	.A(FE_PHN337_n86));
   INVX1 U1674 (.Y(n2388), 
	.A(n879));
   AND2X1 U1675 (.Y(n1396), 
	.B(n1300), 
	.A(FE_OFCN290_n1391));
   INVX1 U1676 (.Y(n2389), 
	.A(n1396));
   AND2X1 U1677 (.Y(n1451), 
	.B(n1312), 
	.A(FE_OFCN289_n1437));
   INVX1 U1678 (.Y(n2390), 
	.A(n1451));
   AND2X1 U1679 (.Y(n1358), 
	.B(DIN[7]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1680 (.Y(n2391), 
	.A(n1358));
   AND2X1 U1681 (.Y(n1381), 
	.B(FE_OFCN319_n1371), 
	.A(mem[89]));
   INVX1 U1682 (.Y(n2392), 
	.A(n1381));
   AND2X1 U1683 (.Y(n1428), 
	.B(n1417), 
	.A(FE_OFCN134_mem_56_));
   INVX1 U1684 (.Y(n2393), 
	.A(n1428));
   AND2X1 U1685 (.Y(n1476), 
	.B(FE_OFCN317_n1463), 
	.A(mem[22]));
   INVX1 U1686 (.Y(n2394), 
	.A(n1476));
   OR2X1 U1688 (.Y(n1095), 
	.B(FE_OFCN38_mem_117_), 
	.A(mem[118]));
   INVX1 U1689 (.Y(n2396), 
	.A(n1095));
   OR2X1 U1691 (.Y(n1159), 
	.B(FE_OFCN118_mem_85_), 
	.A(FE_OFCN117_mem_86_));
   INVX1 U1692 (.Y(n2398), 
	.A(n1159));
   OR2X2 U1694 (.Y(n1288), 
	.B(mem[53]), 
	.A(mem[54]));
   INVX2 U1695 (.Y(n2400), 
	.A(n1288));
   AND2X1 U1701 (.Y(n1506), 
	.B(DIN[3]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1702 (.Y(n2406), 
	.A(n1506));
   AND2X1 U1703 (.Y(n1327), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN41_mem_114_));
   INVX1 U1704 (.Y(n2407), 
	.A(n1327));
   AND2X1 U1705 (.Y(n1393), 
	.B(n251), 
	.A(n1391));
   INVX1 U1706 (.Y(n2408), 
	.A(n1393));
   AND2X1 U1707 (.Y(n1450), 
	.B(n1310), 
	.A(FE_OFCN289_n1437));
   INVX1 U1708 (.Y(n2409), 
	.A(n1450));
   AND2X1 U1709 (.Y(n1363), 
	.B(DIN[4]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1710 (.Y(n2410), 
	.A(n1363));
   AND2X1 U1711 (.Y(n1380), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN113_mem_90_));
   INVX1 U1712 (.Y(n2411), 
	.A(n1380));
   AND2X1 U1713 (.Y(n1427), 
	.B(n1417), 
	.A(mem[57]));
   INVX1 U1714 (.Y(n2412), 
	.A(n1427));
   AND2X1 U1715 (.Y(n1474), 
	.B(FE_OFCN317_n1463), 
	.A(mem[24]));
   INVX1 U1716 (.Y(n2413), 
	.A(n1474));
   AND2X1 U1718 (.Y(n890), 
	.B(n2666), 
	.A(n84));
   INVX1 U1719 (.Y(n2415), 
	.A(n890));
   OR2X2 U1721 (.Y(n1224), 
	.B(mem[22]), 
	.A(mem[23]));
   INVX2 U1722 (.Y(n2417), 
	.A(n1224));
   AND2X1 U1725 (.Y(n1042), 
	.B(n2467), 
	.A(n2501));
   INVX1 U1726 (.Y(n2420), 
	.A(n1042));
   AND2X1 U1727 (.Y(n1041), 
	.B(n2526), 
	.A(n2443));
   INVX1 U1728 (.Y(n2421), 
	.A(n1041));
   AND2X1 U1729 (.Y(n1104), 
	.B(DIN[13]), 
	.A(FE_OFCN38_mem_117_));
   INVX1 U1730 (.Y(n2422), 
	.A(n1104));
   AND2X1 U1731 (.Y(n1168), 
	.B(DIN[13]), 
	.A(mem[85]));
   INVX1 U1732 (.Y(n2423), 
	.A(n1168));
   AND2X1 U1733 (.Y(n1297), 
	.B(DIN[13]), 
	.A(mem[53]));
   INVX2 U1734 (.Y(n2424), 
	.A(n1297));
   OR2X1 U1735 (.Y(n2594), 
	.B(n2595), 
	.A(n1037));
   OR2X1 U1736 (.Y(n2595), 
	.B(n1483), 
	.A(n904));
   AND2X1 U1737 (.Y(n1495), 
	.B(n1306), 
	.A(FE_OFCN288_n1485));
   INVX1 U1738 (.Y(n2425), 
	.A(n1495));
   AND2X1 U1739 (.Y(n1507), 
	.B(DIN[2]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1740 (.Y(n2426), 
	.A(n1507));
   AND2X1 U1741 (.Y(n1329), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN42_mem_113_));
   INVX1 U1742 (.Y(n2427), 
	.A(n1329));
   AND2X1 U1743 (.Y(n1392), 
	.B(n252), 
	.A(n1391));
   INVX1 U1744 (.Y(n2428), 
	.A(n1392));
   AND2X1 U1745 (.Y(n1442), 
	.B(n1300), 
	.A(FE_OFCN289_n1437));
   INVX1 U1746 (.Y(n2429), 
	.A(n1442));
   AND2X1 U1747 (.Y(n1364), 
	.B(DIN[3]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1748 (.Y(n2430), 
	.A(n1364));
   AND2X1 U1749 (.Y(n1384), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN117_mem_86_));
   INVX1 U1750 (.Y(n2431), 
	.A(n1384));
   AND2X1 U1751 (.Y(n1429), 
	.B(FE_OFCN318_n1417), 
	.A(mem[55]));
   INVX1 U1752 (.Y(n2432), 
	.A(n1429));
   AND2X1 U1753 (.Y(n1477), 
	.B(FE_OFCN317_n1463), 
	.A(mem[21]));
   INVX1 U1754 (.Y(n2433), 
	.A(n1477));
   AND2X1 U1755 (.Y(n900), 
	.B(n2666), 
	.A(FE_PHN340_j_3_));
   INVX1 U1756 (.Y(n2434), 
	.A(n900));
   AND2X1 U1758 (.Y(n1105), 
	.B(DIN[14]), 
	.A(FE_OFCN37_mem_118_));
   INVX1 U1759 (.Y(n2436), 
	.A(n1105));
   AND2X1 U1760 (.Y(n1075), 
	.B(DIN[13]), 
	.A(FE_OFCN97_mem_101_));
   INVX1 U1761 (.Y(n2437), 
	.A(n1075));
   AND2X1 U1762 (.Y(n1139), 
	.B(DIN[13]), 
	.A(mem[69]));
   INVX1 U1763 (.Y(n2438), 
	.A(n1139));
   AND2X1 U1764 (.Y(n1233), 
	.B(DIN[15]), 
	.A(mem[23]));
   INVX1 U1765 (.Y(n2439), 
	.A(n1233));
   AND2X1 U1766 (.Y(n1298), 
	.B(DIN[14]), 
	.A(FE_OFCN136_mem_54_));
   INVX2 U1767 (.Y(n2440), 
	.A(n1298));
   AND2X1 U1768 (.Y(n1268), 
	.B(DIN[13]), 
	.A(FE_OFCN71_mem_37_));
   INVX2 U1769 (.Y(n2441), 
	.A(n1268));
   AND2X1 U1770 (.Y(n1277), 
	.B(DIN[10]), 
	.A(FE_OFCN140_mem_50_));
   INVX2 U1771 (.Y(n2442), 
	.A(n1277));
   AND2X1 U1772 (.Y(n948), 
	.B(n1143), 
	.A(n1142));
   INVX1 U1773 (.Y(n2443), 
	.A(n948));
   AND2X1 U1774 (.Y(n1508), 
	.B(DIN[1]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1775 (.Y(n2444), 
	.A(n1508));
   AND2X1 U1776 (.Y(n1305), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN30_mem_125_));
   INVX1 U1777 (.Y(n2445), 
	.A(n1305));
   AND2X1 U1778 (.Y(n1331), 
	.B(FE_OFCN320_n1021), 
	.A(mem[112]));
   INVX1 U1779 (.Y(n2446), 
	.A(n1331));
   AND2X1 U1780 (.Y(n876), 
	.B(n2827), 
	.A(match_addr[2]));
   INVX1 U1781 (.Y(n2447), 
	.A(n876));
   AND2X1 U1782 (.Y(n1403), 
	.B(n1308), 
	.A(n1391));
   INVX1 U1783 (.Y(n2448), 
	.A(n1403));
   AND2X1 U1784 (.Y(n1438), 
	.B(n252), 
	.A(n1437));
   INVX1 U1785 (.Y(n2449), 
	.A(n1438));
   AND2X1 U1786 (.Y(n1365), 
	.B(DIN[2]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1787 (.Y(n2450), 
	.A(n1365));
   AND2X1 U1788 (.Y(n1389), 
	.B(FE_OFCN319_n1371), 
	.A(mem[81]));
   INVX1 U1789 (.Y(n2451), 
	.A(n1389));
   AND2X1 U1790 (.Y(n1430), 
	.B(FE_OFCN318_n1417), 
	.A(FE_OFCN136_mem_54_));
   INVX1 U1791 (.Y(n2452), 
	.A(n1430));
   AND2X1 U1792 (.Y(n1478), 
	.B(FE_OFCN317_n1463), 
	.A(mem[20]));
   INVX1 U1793 (.Y(n2453), 
	.A(n1478));
   AND2X1 U1794 (.Y(n1402), 
	.B(n1306), 
	.A(FE_OFCN290_n1391));
   INVX1 U1795 (.Y(n2454), 
	.A(n1402));
   AND2X1 U1796 (.Y(n1106), 
	.B(DIN[12]), 
	.A(mem[116]));
   INVX1 U1797 (.Y(n2455), 
	.A(n1106));
   AND2X1 U1798 (.Y(n1169), 
	.B(DIN[14]), 
	.A(FE_OFCN117_mem_86_));
   INVX1 U1799 (.Y(n2456), 
	.A(n1169));
   AND2X1 U1800 (.Y(n1140), 
	.B(DIN[14]), 
	.A(FE_OFCN54_mem_70_));
   INVX1 U1801 (.Y(n2457), 
	.A(n1140));
   AND2X2 U1802 (.Y(n1204), 
	.B(DIN[15]), 
	.A(mem[7]));
   INVX1 U1803 (.Y(n2458), 
	.A(n1204));
   AND2X1 U1804 (.Y(n1234), 
	.B(DIN[13]), 
	.A(mem[21]));
   INVX2 U1805 (.Y(n2459), 
	.A(n1234));
   AND2X1 U1806 (.Y(n1269), 
	.B(DIN[14]), 
	.A(mem[38]));
   INVX2 U1807 (.Y(n2460), 
	.A(n1269));
   AND2X1 U1808 (.Y(n1084), 
	.B(DIN[10]), 
	.A(FE_OFCN41_mem_114_));
   INVX1 U1809 (.Y(n2461), 
	.A(n1084));
   AND2X1 U1810 (.Y(n1148), 
	.B(DIN[10]), 
	.A(FE_OFCN121_mem_82_));
   INVX1 U1811 (.Y(n2462), 
	.A(n1148));
   AND2X1 U1812 (.Y(n1229), 
	.B(DIN[10]), 
	.A(mem[18]));
   INVX2 U1813 (.Y(n2463), 
	.A(n1229));
   AND2X1 U1814 (.Y(n1115), 
	.B(DIN[10]), 
	.A(FE_OFCN50_mem_66_));
   INVX1 U1815 (.Y(n2464), 
	.A(n1115));
   AND2X2 U1816 (.Y(n1200), 
	.B(DIN[10]), 
	.A(mem[2]));
   INVX1 U1817 (.Y(n2465), 
	.A(n1200));
   AND2X2 U1818 (.Y(n1244), 
	.B(DIN[10]), 
	.A(mem[34]));
   INVX2 U1819 (.Y(n2466), 
	.A(n1244));
   AND2X1 U1820 (.Y(n932), 
	.B(n1044), 
	.A(n1043));
   INVX1 U1821 (.Y(n2467), 
	.A(n932));
   AND2X2 U1822 (.Y(n979), 
	.B(n1272), 
	.A(n1271));
   INVX1 U1823 (.Y(n2468), 
	.A(n979));
   AND2X1 U1824 (.Y(n1483), 
	.B(n2848), 
	.A(last[0]));
   INVX1 U1825 (.Y(n2469), 
	.A(n1483));
   AND2X1 U1828 (.Y(n1509), 
	.B(DIN[0]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1829 (.Y(n2472), 
	.A(n1509));
   AND2X1 U1830 (.Y(n1317), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN36_mem_119_));
   INVX1 U1831 (.Y(n2473), 
	.A(n1317));
   AND2X1 U1832 (.Y(n1412), 
	.B(DIN[4]), 
	.A(FE_OFCN290_n1391));
   INVX1 U1833 (.Y(n2474), 
	.A(n1412));
   AND2X1 U1834 (.Y(n1449), 
	.B(n1308), 
	.A(FE_OFCN289_n1437));
   INVX1 U1835 (.Y(n2475), 
	.A(n1449));
   AND2X1 U1836 (.Y(n1366), 
	.B(DIN[1]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1837 (.Y(n2476), 
	.A(n1366));
   AND2X1 U1838 (.Y(n1390), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN123_mem_80_));
   INVX1 U1839 (.Y(n2477), 
	.A(n1390));
   AND2X1 U1840 (.Y(n1423), 
	.B(FE_OFCN318_n1417), 
	.A(mem[61]));
   INVX1 U1841 (.Y(n2478), 
	.A(n1423));
   AND2X1 U1842 (.Y(n1434), 
	.B(FE_OFCN318_n1417), 
	.A(FE_OFCN140_mem_50_));
   INVX1 U1843 (.Y(n2479), 
	.A(n1434));
   AND2X2 U1844 (.Y(n1481), 
	.B(n1463), 
	.A(mem[17]));
   INVX1 U1845 (.Y(n2480), 
	.A(n1481));
   AND2X1 U1846 (.Y(n873), 
	.B(n2827), 
	.A(match_addr[1]));
   INVX1 U1847 (.Y(n2481), 
	.A(n873));
   AND2X1 U1848 (.Y(n1492), 
	.B(n1302), 
	.A(FE_OFCN288_n1485));
   INVX1 U1849 (.Y(n2482), 
	.A(n1492));
   AND2X1 U1850 (.Y(n1400), 
	.B(n1304), 
	.A(FE_OFCN290_n1391));
   INVX1 U1851 (.Y(n2483), 
	.A(n1400));
   AND2X1 U1852 (.Y(n1448), 
	.B(n1306), 
	.A(FE_OFCN289_n1437));
   INVX1 U1853 (.Y(n2484), 
	.A(n1448));
   AND2X1 U1854 (.Y(n1076), 
	.B(DIN[14]), 
	.A(FE_OFCN96_mem_102_));
   INVX1 U1855 (.Y(n2485), 
	.A(n1076));
   AND2X1 U1856 (.Y(n1170), 
	.B(DIN[12]), 
	.A(mem[84]));
   INVX1 U1857 (.Y(n2486), 
	.A(n1170));
   AND2X1 U1858 (.Y(n1141), 
	.B(DIN[12]), 
	.A(FE_OFCN52_mem_68_));
   INVX1 U1859 (.Y(n2487), 
	.A(n1141));
   AND2X2 U1860 (.Y(n1206), 
	.B(DIN[14]), 
	.A(mem[6]));
   INVX1 U1861 (.Y(n2488), 
	.A(n1206));
   AND2X2 U1862 (.Y(n1235), 
	.B(DIN[14]), 
	.A(mem[22]));
   INVX2 U1863 (.Y(n2489), 
	.A(n1235));
   AND2X1 U1864 (.Y(n1299), 
	.B(DIN[12]), 
	.A(FE_OFCN138_mem_52_));
   INVX2 U1865 (.Y(n2490), 
	.A(n1299));
   AND2X1 U1866 (.Y(n1270), 
	.B(DIN[12]), 
	.A(mem[36]));
   INVX2 U1867 (.Y(n2491), 
	.A(n1270));
   AND2X1 U1868 (.Y(n1147), 
	.B(DIN[11]), 
	.A(FE_OFCN120_mem_83_));
   INVX1 U1869 (.Y(n2492), 
	.A(n1147));
   AND2X2 U1870 (.Y(n1213), 
	.B(DIN[8]), 
	.A(mem[16]));
   INVX2 U1871 (.Y(n2493), 
	.A(n1213));
   AND2X1 U1872 (.Y(n1276), 
	.B(DIN[11]), 
	.A(mem[51]));
   INVX1 U1873 (.Y(n2494), 
	.A(n1276));
   AND2X1 U1874 (.Y(n1051), 
	.B(DIN[10]), 
	.A(mem[98]));
   INVX1 U1875 (.Y(n2495), 
	.A(n1051));
   AND2X1 U1876 (.Y(n1133), 
	.B(DIN[9]), 
	.A(FE_OFCN49_mem_65_));
   INVX1 U1877 (.Y(n2496), 
	.A(n1133));
   AND2X2 U1878 (.Y(n1178), 
	.B(DIN[12]), 
	.A(FE_OFCN17_mem_4_));
   INVX1 U1879 (.Y(n2497), 
	.A(n1178));
   AND2X2 U1880 (.Y(n1262), 
	.B(DIN[9]), 
	.A(FE_OFCN67_mem_33_));
   INVX1 U1881 (.Y(n2498), 
	.A(n1262));
   AND2X1 U1884 (.Y(n914), 
	.B(n1079), 
	.A(n1078));
   INVX1 U1885 (.Y(n2501), 
	.A(n914));
   AND2X1 U1886 (.Y(n887), 
	.B(n906), 
	.A(FE_OFCN255_n897));
   INVX1 U1887 (.Y(n2502), 
	.A(n887));
   AND2X1 U1890 (.Y(n1321), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN38_mem_117_));
   INVX1 U1891 (.Y(n2505), 
	.A(n1321));
   AND2X1 U1892 (.Y(n1367), 
	.B(DIN[0]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1893 (.Y(n2506), 
	.A(n1367));
   AND2X1 U1894 (.Y(n1377), 
	.B(FE_OFCN319_n1371), 
	.A(mem[93]));
   INVX1 U1895 (.Y(n2507), 
	.A(n1377));
   AND2X1 U1896 (.Y(n1388), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN121_mem_82_));
   INVX1 U1897 (.Y(n2508), 
	.A(n1388));
   AND2X1 U1898 (.Y(n1435), 
	.B(n1417), 
	.A(mem[49]));
   INVX1 U1899 (.Y(n2509), 
	.A(n1435));
   AND2X1 U1900 (.Y(n1468), 
	.B(FE_OFCN317_n1463), 
	.A(mem[30]));
   INVX1 U1901 (.Y(n2510), 
	.A(n1468));
   AND2X1 U1902 (.Y(n1479), 
	.B(n1463), 
	.A(mem[19]));
   INVX1 U1903 (.Y(n2511), 
	.A(n1479));
   AND2X1 U1904 (.Y(n870), 
	.B(n2827), 
	.A(match_addr[0]));
   INVX1 U1905 (.Y(n2512), 
	.A(n870));
   AND2X1 U1906 (.Y(n1490), 
	.B(n1300), 
	.A(FE_OFCN288_n1485));
   INVX1 U1907 (.Y(n2513), 
	.A(n1490));
   AND2X1 U1908 (.Y(n1395), 
	.B(n250), 
	.A(n1391));
   INVX1 U1909 (.Y(n2514), 
	.A(n1395));
   AND2X1 U1910 (.Y(n1455), 
	.B(DIN[6]), 
	.A(FE_OFCN289_n1437));
   INVX1 U1911 (.Y(n2515), 
	.A(n1455));
   AND2X1 U1912 (.Y(n1446), 
	.B(n1304), 
	.A(FE_OFCN289_n1437));
   INVX1 U1913 (.Y(n2516), 
	.A(n1446));
   AND2X1 U1914 (.Y(n1342), 
	.B(n1302), 
	.A(FE_OFCN291_n1335));
   INVX1 U1915 (.Y(n2517), 
	.A(n1342));
   AND2X1 U1916 (.Y(n1077), 
	.B(DIN[12]), 
	.A(FE_OFCN98_mem_100_));
   INVX1 U1917 (.Y(n2518), 
	.A(n1077));
   AND2X1 U1918 (.Y(n1205), 
	.B(DIN[13]), 
	.A(mem[5]));
   INVX2 U1919 (.Y(n2519), 
	.A(n1205));
   AND2X1 U1920 (.Y(n1100), 
	.B(DIN[8]), 
	.A(FE_OFCN43_mem_112_));
   INVX1 U1921 (.Y(n2520), 
	.A(n1100));
   AND2X1 U1922 (.Y(n1164), 
	.B(DIN[8]), 
	.A(FE_OFCN123_mem_80_));
   INVX1 U1923 (.Y(n2521), 
	.A(n1164));
   AND2X1 U1924 (.Y(n1293), 
	.B(DIN[8]), 
	.A(mem[48]));
   INVX2 U1925 (.Y(n2522), 
	.A(n1293));
   AND2X1 U1926 (.Y(n1228), 
	.B(DIN[9]), 
	.A(mem[17]));
   INVX2 U1927 (.Y(n2523), 
	.A(n1228));
   AND2X1 U1928 (.Y(n1069), 
	.B(DIN[9]), 
	.A(mem[97]));
   INVX1 U1929 (.Y(n2524), 
	.A(n1069));
   AND2X1 U1931 (.Y(n964), 
	.B(n1108), 
	.A(n1107));
   INVX1 U1932 (.Y(n2526), 
	.A(n964));
   AND2X2 U1933 (.Y(n995), 
	.B(n1237), 
	.A(n1236));
   INVX1 U1934 (.Y(n2527), 
	.A(n995));
   OR2X1 U1935 (.Y(n885), 
	.B(n2798), 
	.A(n2800));
   INVX1 U1936 (.Y(n2528), 
	.A(n885));
   INVX1 U1945 (.Y(n2537), 
	.A(FE_PSN328_n1003));
   AND2X1 U1953 (.Y(n1319), 
	.B(FE_OFCN320_n1021), 
	.A(FE_OFCN37_mem_118_));
   INVX1 U1954 (.Y(n2545), 
	.A(n1319));
   AND2X1 U1955 (.Y(n1385), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN118_mem_85_));
   INVX1 U1956 (.Y(n2546), 
	.A(n1385));
   AND2X1 U1957 (.Y(n1436), 
	.B(FE_OFCN318_n1417), 
	.A(mem[48]));
   INVX1 U1958 (.Y(n2547), 
	.A(n1436));
   AND2X1 U1959 (.Y(n1469), 
	.B(FE_OFCN317_n1463), 
	.A(mem[29]));
   INVX1 U1960 (.Y(n2548), 
	.A(n1469));
   AND2X2 U1961 (.Y(n1480), 
	.B(n1463), 
	.A(mem[18]));
   INVX1 U1962 (.Y(n2549), 
	.A(n1480));
   AND2X1 U1963 (.Y(n1501), 
	.B(DIN[7]), 
	.A(FE_OFCN288_n1485));
   INVX1 U1964 (.Y(n2550), 
	.A(n1501));
   AND2X1 U1965 (.Y(n1409), 
	.B(DIN[6]), 
	.A(FE_OFCN290_n1391));
   INVX1 U1966 (.Y(n2551), 
	.A(n1409));
   AND2X1 U1967 (.Y(n1398), 
	.B(n1302), 
	.A(FE_OFCN290_n1391));
   INVX1 U1968 (.Y(n2552), 
	.A(n1398));
   AND2X1 U1969 (.Y(n1441), 
	.B(n250), 
	.A(n1437));
   INVX1 U1970 (.Y(n2553), 
	.A(n1441));
   AND2X1 U1971 (.Y(n1345), 
	.B(n1304), 
	.A(FE_OFCN291_n1335));
   INVX1 U1972 (.Y(n2554), 
	.A(n1345));
   AND2X1 U1973 (.Y(n1360), 
	.B(DIN[6]), 
	.A(FE_OFCN291_n1335));
   INVX1 U1974 (.Y(n2555), 
	.A(n1360));
   INVX1 U1975 (.Y(n2556), 
	.A(n1781));
   INVX1 U1976 (.Y(n2557), 
	.A(n874));
   INVX1 U1977 (.Y(n2558), 
	.A(n2984));
   AND2X1 U1978 (.Y(n2984), 
	.B(n2622), 
	.A(n2699));
   INVX1 U1979 (.Y(n2559), 
	.A(n1083));
   AND2X1 U1980 (.Y(n1071), 
	.B(DIN[8]), 
	.A(mem[96]));
   INVX1 U1981 (.Y(n2560), 
	.A(n1071));
   AND2X1 U1982 (.Y(n1135), 
	.B(DIN[8]), 
	.A(FE_OFCN48_mem_64_));
   INVX1 U1983 (.Y(n2561), 
	.A(n1135));
   AND2X2 U1984 (.Y(n1180), 
	.B(DIN[8]), 
	.A(FE_OFCN21_mem_0_));
   INVX1 U1985 (.Y(n2562), 
	.A(n1180));
   AND2X2 U1986 (.Y(n1264), 
	.B(DIN[8]), 
	.A(mem[32]));
   INVX2 U1987 (.Y(n2563), 
	.A(n1264));
   AND2X1 U1988 (.Y(n1648), 
	.B(n2774), 
	.A(rank[8]));
   INVX1 U1989 (.Y(n2564), 
	.A(n1648));
   AND2X1 U2011 (.Y(n976), 
	.B(n967), 
	.A(n2809));
   INVX2 U2012 (.Y(n2586), 
	.A(n976));
   AND2X1 U2018 (.Y(n1009), 
	.B(n2961), 
	.A(n998));
   INVX2 U2019 (.Y(n2592), 
	.A(n1009));
   AND2X2 U2020 (.Y(n998), 
	.B(n1003), 
	.A(FE_OFCN3_matchN_2_));
   AND2X1 U2024 (.Y(n945), 
	.B(n936), 
	.A(n2805));
   INVX2 U2025 (.Y(n2598), 
	.A(n945));
   AND2X1 U2026 (.Y(n1027), 
	.B(n1021), 
	.A(matchN[21]));
   INVX1 U2027 (.Y(n2599), 
	.A(n1027));
   AND2X1 U2028 (.Y(n1383), 
	.B(FE_OFCN319_n1371), 
	.A(FE_OFCN116_mem_87_));
   INVX1 U2029 (.Y(n2600), 
	.A(n1383));
   AND2X1 U2030 (.Y(n1431), 
	.B(FE_OFCN318_n1417), 
	.A(mem[53]));
   INVX1 U2031 (.Y(n2601), 
	.A(n1431));
   AND2X2 U2032 (.Y(n1482), 
	.B(n1463), 
	.A(mem[16]));
   INVX1 U2033 (.Y(n2602), 
	.A(n1482));
   AND2X1 U2034 (.Y(n1494), 
	.B(n1304), 
	.A(FE_OFCN288_n1485));
   INVX1 U2035 (.Y(n2603), 
	.A(n1494));
   AND2X1 U2036 (.Y(n1503), 
	.B(DIN[6]), 
	.A(FE_OFCN288_n1485));
   INVX1 U2037 (.Y(n2604), 
	.A(n1503));
   AND2X1 U2038 (.Y(n1411), 
	.B(DIN[5]), 
	.A(FE_OFCN290_n1391));
   INVX1 U2039 (.Y(n2605), 
	.A(n1411));
   AND2X1 U2040 (.Y(n1457), 
	.B(DIN[5]), 
	.A(FE_OFCN289_n1437));
   INVX1 U2041 (.Y(n2606), 
	.A(n1457));
   AND2X1 U2042 (.Y(n1444), 
	.B(n1302), 
	.A(FE_OFCN289_n1437));
   INVX1 U2043 (.Y(n2607), 
	.A(n1444));
   AND2X1 U2044 (.Y(n1348), 
	.B(n1306), 
	.A(FE_OFCN291_n1335));
   INVX1 U2045 (.Y(n2608), 
	.A(n1348));
   AND2X1 U2046 (.Y(n1362), 
	.B(DIN[5]), 
	.A(FE_OFCN291_n1335));
   INVX1 U2047 (.Y(n2609), 
	.A(n1362));
   BUFX2 U2048 (.Y(match_addr[2]), 
	.A(FE_OFCN44_n3000));
   BUFX2 U2049 (.Y(match_addr[1]), 
	.A(FE_OFCN168_n3001));
   BUFX2 U2050 (.Y(match_addr[0]), 
	.A(FE_OFCN175_n3002));
   AND2X1 U2051 (.Y(n1049), 
	.B(DIN[11]), 
	.A(FE_OFCN99_mem_99_));
   INVX1 U2052 (.Y(n2613), 
	.A(n1049));
   AND2X1 U2053 (.Y(n1113), 
	.B(DIN[11]), 
	.A(mem[67]));
   INVX1 U2054 (.Y(n2614), 
	.A(n1113));
   AND2X1 U2055 (.Y(n1242), 
	.B(DIN[11]), 
	.A(mem[35]));
   INVX1 U2056 (.Y(n2615), 
	.A(n1242));
   AND2X2 U2057 (.Y(n1198), 
	.B(DIN[9]), 
	.A(mem[1]));
   INVX1 U2058 (.Y(n2616), 
	.A(n1198));
   AND2X1 U2064 (.Y(n2986), 
	.B(n2823), 
	.A(n236));
   INVX1 U2065 (.Y(n2622), 
	.A(n2986));
   AND2X1 U2109 (.Y(n880), 
	.B(n901), 
	.A(n2796));
   INVX4 U2110 (.Y(n2666), 
	.A(n880));
   INVX1 U2111 (.Y(n2667), 
	.A(n905));
   AND2X1 U2112 (.Y(n1439), 
	.B(n251), 
	.A(n1437));
   INVX1 U2113 (.Y(n2668), 
	.A(n1439));
   AND2X1 U2114 (.Y(n1338), 
	.B(n250), 
	.A(FE_OFCN291_n1335));
   INVX1 U2115 (.Y(n2669), 
	.A(n1338));
   INVX1 U2116 (.Y(n2670), 
	.A(n1099));
   INVX1 U2117 (.Y(n2671), 
	.A(n1163));
   INVX1 U2118 (.Y(n2672), 
	.A(n1212));
   INVX1 U2119 (.Y(n2673), 
	.A(n1292));
   AND2X1 U2145 (.Y(n2985), 
	.B(n2988), 
	.A(n2987));
   INVX1 U2146 (.Y(n2699), 
	.A(n2985));
   AND2X1 U2177 (.Y(n903), 
	.B(n2946), 
	.A(EN));
   INVX1 U2178 (.Y(n2730), 
	.A(n903));
   AND2X1 U2187 (.Y(n1308), 
	.B(DIN[11]), 
	.A(DIN[3]));
   INVX1 U2188 (.Y(n2739), 
	.A(n1308));
   AND2X1 U2189 (.Y(n1310), 
	.B(DIN[10]), 
	.A(DIN[2]));
   INVX1 U2190 (.Y(n2740), 
	.A(n1310));
   AND2X1 U2191 (.Y(n1312), 
	.B(DIN[9]), 
	.A(DIN[1]));
   INVX1 U2192 (.Y(n2741), 
	.A(n1312));
   AND2X1 U2193 (.Y(n1314), 
	.B(DIN[8]), 
	.A(DIN[0]));
   INVX1 U2194 (.Y(n2742), 
	.A(n1314));
   AND2X1 U2195 (.Y(n1300), 
	.B(DIN[15]), 
	.A(DIN[7]));
   INVX1 U2196 (.Y(n2743), 
	.A(n1300));
   AND2X1 U2197 (.Y(n1306), 
	.B(DIN[12]), 
	.A(DIN[4]));
   INVX1 U2198 (.Y(n2744), 
	.A(n1306));
   AND2X1 U2199 (.Y(n1302), 
	.B(DIN[14]), 
	.A(DIN[6]));
   INVX1 U2200 (.Y(n2745), 
	.A(n1302));
   AND2X1 U2201 (.Y(n1304), 
	.B(DIN[13]), 
	.A(DIN[5]));
   INVX1 U2202 (.Y(n2746), 
	.A(n1304));
   AND2X1 U2205 (.Y(n929), 
	.B(n2802), 
	.A(n2803));
   INVX2 U2206 (.Y(n2749), 
	.A(n929));
   AND2X1 U2208 (.Y(n992), 
	.B(n2811), 
	.A(n2810));
   INVX2 U2209 (.Y(n2751), 
	.A(n992));
   INVX1 U2210 (.Y(n2752), 
	.A(n868));
   AND2X1 U2212 (.Y(n961), 
	.B(n2806), 
	.A(n2807));
   INVX2 U2213 (.Y(n2754), 
	.A(n961));
   INVX1 U2214 (.Y(n2813), 
	.A(n251));
   INVX1 U2215 (.Y(n2814), 
	.A(n252));
   INVX1 U2219 (.Y(n2790), 
	.A(reset));
   INVX1 U2220 (.Y(n2789), 
	.A(reset));
   INVX1 U2221 (.Y(n2788), 
	.A(reset));
   INVX1 U2222 (.Y(n2787), 
	.A(reset));
   INVX1 U2223 (.Y(n2785), 
	.A(reset));
   INVX1 U2224 (.Y(n2786), 
	.A(reset));
   INVX1 U2225 (.Y(n2784), 
	.A(reset));
   INVX1 U2226 (.Y(n2783), 
	.A(reset));
   INVX1 U2227 (.Y(n2782), 
	.A(reset));
   INVX1 U2228 (.Y(n2781), 
	.A(reset));
   INVX1 U2229 (.Y(n2780), 
	.A(reset));
   INVX1 U2230 (.Y(n2779), 
	.A(reset));
   INVX4 U2231 (.Y(n2804), 
	.A(FE_OFCN263_n886));
   INVX2 U2232 (.Y(n2800), 
	.A(FE_OFCN268_n892));
   INVX2 U2233 (.Y(n2808), 
	.A(n906));
   INVX1 U2234 (.Y(n2801), 
	.A(FE_PSN331_FE_OFCN261_n888));
   INVX1 U2235 (.Y(n2816), 
	.A(n250));
   INVX1 U2236 (.Y(n2832), 
	.A(n1660));
   INVX1 U2237 (.Y(n2836), 
	.A(n1617));
   INVX1 U2238 (.Y(n2834), 
	.A(n1639));
   INVX1 U2239 (.Y(n2838), 
	.A(n1596));
   INVX1 U2240 (.Y(n2830), 
	.A(n1534));
   INVX1 U2241 (.Y(n2840), 
	.A(n1575));
   INVX1 U2242 (.Y(n2842), 
	.A(n1548));
   INVX1 U2243 (.Y(n2828), 
	.A(n1681));
   INVX1 U2247 (.Y(n2873), 
	.A(n1037));
   INVX1 U2248 (.Y(n2812), 
	.A(FE_OFCN250_n1005));
   OR2X2 U2249 (.Y(n916), 
	.B(n912), 
	.A(FE_PHN336_n2878));
   INVX1 U2250 (.Y(n2802), 
	.A(FE_OFCN267_n928));
   INVX2 U2251 (.Y(n2806), 
	.A(n952));
   INVX2 U2252 (.Y(n2811), 
	.A(n983));
   INVX1 U2253 (.Y(n2798), 
	.A(n908));
   AND2X1 U2254 (.Y(n1017), 
	.B(n1173), 
	.A(n1172));
   AND2X1 U2255 (.Y(n2987), 
	.B(n233), 
	.A(n235));
   INVX1 U2257 (.Y(n2874), 
	.A(FE_OFCN183_n1522));
   INVX1 U2258 (.Y(n2846), 
	.A(FE_OFCN229_n1368));
   INVX1 U2259 (.Y(n2847), 
	.A(FE_OFCN228_n1369));
   INVX2 U2260 (.Y(n2961), 
	.A(matchN[5]));
   INVX1 U2261 (.Y(n2962), 
	.A(matchN[4]));
   INVX2 U2262 (.Y(n2966), 
	.A(mem[19]));
   AND2X2 U2263 (.Y(n1183), 
	.B(n2859), 
	.A(DIN[11]));
   INVX2 U2264 (.Y(n2805), 
	.A(n953));
   INVX1 U2265 (.Y(n2797), 
	.A(n881));
   INVX2 U2266 (.Y(n2809), 
	.A(n984));
   OR2X2 U2267 (.Y(n917), 
	.B(n919), 
	.A(n2879));
   INVX2 U2268 (.Y(n2799), 
	.A(n921));
   INVX2 U2269 (.Y(n2810), 
	.A(n999));
   INVX1 U2270 (.Y(n2807), 
	.A(n968));
   INVX1 U2271 (.Y(n2803), 
	.A(n937));
   AND2X2 U2272 (.Y(n1011), 
	.B(n1208), 
	.A(n1207));
   AND2X2 U2273 (.Y(n1216), 
	.B(n2963), 
	.A(DIN[11]));
   INVX1 U2274 (.Y(n2795), 
	.A(FE_PHN334_FE_OFCN322_n882));
   AND2X2 U2275 (.Y(n1247), 
	.B(n2924), 
	.A(DIN[15]));
   INVX2 U2276 (.Y(n2957), 
	.A(FE_OFCN135_mem_55_));
   INVX1 U2277 (.Y(n2950), 
	.A(mem[87]));
   AND2X1 U2278 (.Y(n1118), 
	.B(n2905), 
	.A(DIN[15]));
   INVX2 U2279 (.Y(n2964), 
	.A(mem[21]));
   INVX2 U2280 (.Y(n2965), 
	.A(mem[20]));
   INVX2 U2281 (.Y(n2853), 
	.A(FE_OFCN4_matchN_1_));
   INVX4 U2282 (.Y(n2854), 
	.A(matchN[0]));
   INVX2 U2283 (.Y(n2967), 
	.A(n1221));
   INVX2 U2284 (.Y(n2924), 
	.A(mem[47]));
   INVX2 U2285 (.Y(n2859), 
	.A(mem[11]));
   INVX2 U2286 (.Y(n2867), 
	.A(mem[3]));
   INVX2 U2287 (.Y(n2963), 
	.A(mem[27]));
   INVX1 U2288 (.Y(n2909), 
	.A(mem[32]));
   INVX2 U2289 (.Y(n2870), 
	.A(mem[0]));
   INVX2 U2290 (.Y(n2913), 
	.A(mem[36]));
   INVX1 U2291 (.Y(n2911), 
	.A(mem[34]));
   INVX2 U2292 (.Y(n2865), 
	.A(mem[5]));
   INVX2 U2293 (.Y(n2868), 
	.A(mem[2]));
   INVX2 U2294 (.Y(n2912), 
	.A(mem[35]));
   INVX2 U2295 (.Y(n2910), 
	.A(mem[33]));
   INVX2 U2296 (.Y(n2866), 
	.A(mem[4]));
   INVX2 U2297 (.Y(n2869), 
	.A(mem[1]));
   INVX2 U2298 (.Y(n2852), 
	.A(matchN[2]));
   INVX2 U2299 (.Y(n2862), 
	.A(mem[8]));
   INVX2 U2300 (.Y(n2858), 
	.A(mem[12]));
   INVX2 U2301 (.Y(n2860), 
	.A(mem[10]));
   INVX2 U2302 (.Y(n2861), 
	.A(mem[9]));
   AND2X2 U2303 (.Y(n1280), 
	.B(n2956), 
	.A(DIN[15]));
   AND2X1 U2304 (.Y(n1151), 
	.B(n2949), 
	.A(DIN[15]));
   AND2X1 U2305 (.Y(n1054), 
	.B(n2930), 
	.A(DIN[15]));
   INVX1 U2306 (.Y(n2881), 
	.A(FE_OFCN36_mem_119_));
   INVX1 U2307 (.Y(n2864), 
	.A(mem[6]));
   INVX1 U2308 (.Y(n2863), 
	.A(mem[7]));
   INVX1 U2309 (.Y(n2857), 
	.A(mem[13]));
   INVX1 U2310 (.Y(n2856), 
	.A(mem[14]));
   INVX1 U2311 (.Y(n2855), 
	.A(mem[15]));
   INVX1 U2312 (.Y(n2915), 
	.A(mem[38]));
   INVX1 U2313 (.Y(n2914), 
	.A(FE_OFCN71_mem_37_));
   INVX1 U2314 (.Y(n2896), 
	.A(mem[70]));
   INVX1 U2315 (.Y(n2895), 
	.A(FE_OFCN53_mem_69_));
   INVX1 U2316 (.Y(n2940), 
	.A(mem[101]));
   INVX1 U2317 (.Y(n2939), 
	.A(FE_OFCN96_mem_102_));
   INVX1 U2318 (.Y(n2925), 
	.A(matchN[6]));
   INVX1 U2319 (.Y(n2923), 
	.A(FE_OFCN80_mem_46_));
   INVX1 U2320 (.Y(n2922), 
	.A(mem[45]));
   INVX1 U2321 (.Y(n2921), 
	.A(mem[44]));
   INVX1 U2322 (.Y(n2906), 
	.A(matchN[12]));
   INVX1 U2323 (.Y(n2904), 
	.A(FE_OFCN61_mem_78_));
   INVX1 U2324 (.Y(n2903), 
	.A(mem[77]));
   INVX1 U2325 (.Y(n2902), 
	.A(mem[76]));
   INVX1 U2326 (.Y(n2933), 
	.A(mem[108]));
   INVX1 U2327 (.Y(n2932), 
	.A(FE_OFCN90_mem_109_));
   INVX1 U2328 (.Y(n2931), 
	.A(mem[110]));
   INVX1 U2329 (.Y(n2833), 
	.A(n1657));
   INVX1 U2330 (.Y(n2837), 
	.A(n1614));
   INVX1 U2331 (.Y(n2835), 
	.A(n1636));
   INVX1 U2332 (.Y(n2839), 
	.A(n1593));
   INVX1 U2333 (.Y(n2831), 
	.A(n1533));
   INVX1 U2334 (.Y(n2841), 
	.A(n1572));
   INVX1 U2335 (.Y(n2843), 
	.A(n1545));
   INVX1 U2336 (.Y(n2829), 
	.A(n1678));
   INVX2 U2337 (.Y(n2958), 
	.A(FE_OFCN138_mem_52_));
   INVX2 U2338 (.Y(n2959), 
	.A(mem[51]));
   INVX1 U2339 (.Y(n2951), 
	.A(FE_OFCN119_mem_84_));
   INVX1 U2340 (.Y(n2952), 
	.A(mem[83]));
   INVX1 U2341 (.Y(n2889), 
	.A(FE_PHN341_last_1_));
   INVX1 U2342 (.Y(n2877), 
	.A(last[2]));
   INVX1 U2343 (.Y(n2851), 
	.A(last[0]));
   INVX2 U2344 (.Y(n2960), 
	.A(n1285));
   INVX1 U2345 (.Y(n2953), 
	.A(n1156));
   INVX4 U2346 (.Y(n2926), 
	.A(matchN[7]));
   INVX1 U2347 (.Y(n2907), 
	.A(FE_OFCN64_matchN_13_));
   INVX1 U2348 (.Y(n2815), 
	.A(FE_OFCN277_n2990));
   AND2X1 U2349 (.Y(n2992), 
	.B(n238), 
	.A(DIN[4]));
   INVX1 U2350 (.Y(n2818), 
	.A(FE_OFCN278_n2993));
   AND2X1 U2351 (.Y(n2995), 
	.B(DIN[5]), 
	.A(DIN[6]));
   INVX1 U2352 (.Y(n2823), 
	.A(FE_OFCN279_n2996));
   AND2X1 U2353 (.Y(n2998), 
	.B(DIN[2]), 
	.A(DIN[1]));
   INVX1 U2354 (.Y(n2955), 
	.A(matchN[10]));
   INVX1 U2355 (.Y(n2948), 
	.A(matchN[16]));
   INVX1 U2356 (.Y(n2905), 
	.A(FE_OFCN62_mem_79_));
   INVX1 U2357 (.Y(n2916), 
	.A(mem[39]));
   INVX1 U2358 (.Y(n2897), 
	.A(FE_OFCN55_mem_71_));
   INVX1 U2359 (.Y(n2954), 
	.A(FE_OFCN124_matchN_11_));
   INVX1 U2360 (.Y(n2947), 
	.A(FE_OFCN105_matchN_17_));
   INVX2 U2361 (.Y(n2956), 
	.A(mem[63]));
   INVX1 U2362 (.Y(n2949), 
	.A(FE_OFCN108_mem_95_));
   INVX1 U2363 (.Y(n2890), 
	.A(mem[64]));
   INVX1 U2364 (.Y(n2894), 
	.A(FE_OFCN52_mem_68_));
   INVX1 U2365 (.Y(n2892), 
	.A(mem[66]));
   INVX1 U2366 (.Y(n2893), 
	.A(FE_OFCN51_mem_67_));
   INVX1 U2367 (.Y(n2891), 
	.A(FE_OFCN49_mem_65_));
   INVX1 U2368 (.Y(n2826), 
	.A(DIN[0]));
   INVX1 U2369 (.Y(n2825), 
	.A(DIN[1]));
   INVX1 U2370 (.Y(n2824), 
	.A(DIN[2]));
   INVX1 U2371 (.Y(n2822), 
	.A(DIN[3]));
   INVX1 U2372 (.Y(n2821), 
	.A(DIN[4]));
   INVX1 U2373 (.Y(n2820), 
	.A(DIN[5]));
   INVX1 U2374 (.Y(n2819), 
	.A(DIN[6]));
   INVX1 U2375 (.Y(n2817), 
	.A(DIN[7]));
   INVX2 U2376 (.Y(n2917), 
	.A(mem[40]));
   INVX2 U2377 (.Y(n2918), 
	.A(mem[41]));
   INVX2 U2378 (.Y(n2919), 
	.A(mem[42]));
   INVX2 U2379 (.Y(n2920), 
	.A(mem[43]));
   INVX1 U2380 (.Y(n2898), 
	.A(FE_OFCN56_mem_72_));
   INVX1 U2381 (.Y(n2899), 
	.A(FE_OFCN57_mem_73_));
   INVX1 U2382 (.Y(n2900), 
	.A(mem[74]));
   INVX1 U2383 (.Y(n2901), 
	.A(FE_OFCN58_mem_75_));
   INVX2 U2384 (.Y(n2927), 
	.A(matchN[8]));
   INVX1 U2385 (.Y(n2908), 
	.A(FE_OFCN65_matchN_14_));
   AND2X1 U2386 (.Y(n1087), 
	.B(n2880), 
	.A(DIN[15]));
   INVX1 U2388 (.Y(n2796), 
	.A(reset));
   INVX1 U2389 (.Y(n2827), 
	.A(EN));
   INVX1 U2390 (.Y(n2844), 
	.A(WE));
   INVX1 U2391 (.Y(n2871), 
	.A(n84));
   INVX1 U2392 (.Y(n88), 
	.A(n2773));
   INVX1 U2393 (.Y(n2884), 
	.A(n1092));
   INVX1 U2394 (.Y(n2968), 
	.A(n85));
   INVX1 U2395 (.Y(n2882), 
	.A(FE_OFCN39_mem_116_));
   INVX1 U2396 (.Y(n2883), 
	.A(mem[115]));
   INVX1 U2397 (.Y(n87), 
	.A(n2774));
   INVX1 U2398 (.Y(n2983), 
	.A(rank[4]));
   INVX1 U2399 (.Y(n2980), 
	.A(rank[10]));
   INVX1 U2400 (.Y(n2977), 
	.A(rank[7]));
   INVX1 U2401 (.Y(n2974), 
	.A(rank[13]));
   INVX1 U2402 (.Y(n2969), 
	.A(rank[22]));
   INVX1 U2403 (.Y(n2888), 
	.A(FE_OFCN47_rank_16_));
   INVX1 U2404 (.Y(n2876), 
	.A(rank[19]));
   INVX1 U2405 (.Y(n2849), 
	.A(rank[1]));
   INVX1 U2406 (.Y(n2982), 
	.A(FE_OFCN177_rank_3_));
   INVX1 U2407 (.Y(n2979), 
	.A(rank[9]));
   INVX1 U2408 (.Y(n2976), 
	.A(rank[6]));
   INVX1 U2409 (.Y(n2973), 
	.A(FE_OFCN166_rank_12_));
   INVX1 U2410 (.Y(n2970), 
	.A(rank[21]));
   INVX1 U2411 (.Y(n2887), 
	.A(FE_OFCN46_rank_15_));
   INVX1 U2412 (.Y(n2875), 
	.A(FE_OFCN23_rank_18_));
   INVX1 U2413 (.Y(n2845), 
	.A(FE_OFCN0_rank_0_));
   INVX1 U2414 (.Y(n2946), 
	.A(FE_OFCN103_m));
   INVX1 U2415 (.Y(n2981), 
	.A(rank[5]));
   INVX1 U2416 (.Y(n2978), 
	.A(rank[11]));
   INVX1 U2417 (.Y(n2975), 
	.A(rank[8]));
   INVX1 U2418 (.Y(n2972), 
	.A(rank[14]));
   INVX1 U2419 (.Y(n2971), 
	.A(rank[23]));
   INVX1 U2420 (.Y(n2886), 
	.A(rank[17]));
   INVX1 U2421 (.Y(n2872), 
	.A(FE_OFCN22_rank_20_));
   INVX1 U2422 (.Y(n2850), 
	.A(rank[2]));
   INVX1 U2423 (.Y(n2885), 
	.A(n86));
   INVX1 U2424 (.Y(n2848), 
	.A(FE_OFCN227_n1525));
   INVX1 U2425 (.Y(n2929), 
	.A(FE_OFCN86_matchN_19_));
   INVX1 U2426 (.Y(n2930), 
	.A(FE_OFCN88_mem_111_));
   INVX1 U2427 (.Y(n2938), 
	.A(FE_OFCN95_mem_103_));
   INVX1 U2428 (.Y(n2880), 
	.A(FE_OFCN28_mem_127_));
   INVX1 U2429 (.Y(n2945), 
	.A(FE_OFCN102_mem_96_));
   INVX1 U2430 (.Y(n2941), 
	.A(mem[100]));
   INVX1 U2431 (.Y(n2943), 
	.A(FE_OFCN100_mem_98_));
   INVX1 U2432 (.Y(n2942), 
	.A(FE_OFCN99_mem_99_));
   INVX1 U2433 (.Y(n2944), 
	.A(FE_OFCN101_mem_97_));
   INVX1 U2434 (.Y(FE_PHN335_n2879), 
	.A(matchN[22]));
   INVX1 U2435 (.Y(n2878), 
	.A(matchN[23]));
   INVX1 U2436 (.Y(n2937), 
	.A(FE_OFCN94_mem_104_));
   INVX1 U2437 (.Y(n2936), 
	.A(mem[105]));
   INVX1 U2438 (.Y(n2935), 
	.A(FE_OFCN93_mem_106_));
   INVX1 U2439 (.Y(n2934), 
	.A(FE_OFCN92_mem_107_));
   INVX1 U2440 (.Y(n2928), 
	.A(FE_OFCN85_matchN_20_));
   MUX2X1 U2441 (.Y(n2755), 
	.S(n85), 
	.B(n2756), 
	.A(n2757));
   MUX2X1 U2442 (.Y(n2758), 
	.S(n85), 
	.B(n2759), 
	.A(n2760));
   MUX2X1 U2443 (.Y(n2761), 
	.S(n85), 
	.B(n2762), 
	.A(n2763));
   MUX2X1 U2444 (.Y(n2764), 
	.S(n85), 
	.B(n2765), 
	.A(n2766));
   MUX2X1 U2445 (.Y(n2767), 
	.S(n85), 
	.B(n2768), 
	.A(n2769));
   MUX2X1 U2446 (.Y(n2770), 
	.S(n85), 
	.B(n2771), 
	.A(n2772));
   MUX2X1 U2447 (.Y(n2757), 
	.S(n84), 
	.B(FE_OFCN23_rank_18_), 
	.A(rank[21]));
   MUX2X1 U2448 (.Y(n2756), 
	.S(n84), 
	.B(FE_OFCN166_rank_12_), 
	.A(FE_OFCN46_rank_15_));
   MUX2X1 U2449 (.Y(n2760), 
	.S(n84), 
	.B(rank[6]), 
	.A(rank[9]));
   MUX2X1 U2450 (.Y(n2759), 
	.S(n84), 
	.B(FE_OFCN0_rank_0_), 
	.A(FE_OFCN177_rank_3_));
   MUX2X1 U2451 (.Y(n89), 
	.S(n86), 
	.B(n2758), 
	.A(n2755));
   MUX2X1 U2452 (.Y(n2763), 
	.S(n84), 
	.B(rank[19]), 
	.A(FE_OFCN162_rank_22_));
   MUX2X1 U2453 (.Y(n2762), 
	.S(n84), 
	.B(FE_OFCN167_rank_13_), 
	.A(FE_OFCN47_rank_16_));
   MUX2X1 U2454 (.Y(n2766), 
	.S(n84), 
	.B(rank[7]), 
	.A(rank[10]));
   MUX2X1 U2455 (.Y(n2765), 
	.S(n84), 
	.B(FE_OFCN1_rank_1_), 
	.A(FE_OFCN178_rank_4_));
   MUX2X1 U2456 (.Y(n2773), 
	.S(n86), 
	.B(n2764), 
	.A(n2761));
   MUX2X1 U2457 (.Y(n2769), 
	.S(n84), 
	.B(FE_OFCN22_rank_20_), 
	.A(FE_OFCN164_rank_23_));
   MUX2X1 U2458 (.Y(n2768), 
	.S(n84), 
	.B(rank[14]), 
	.A(rank[17]));
   MUX2X1 U2459 (.Y(n2772), 
	.S(n84), 
	.B(rank[8]), 
	.A(rank[11]));
   MUX2X1 U2460 (.Y(n2771), 
	.S(n84), 
	.B(FE_OFCN2_rank_2_), 
	.A(rank[5]));
   MUX2X1 U2461 (.Y(n2774), 
	.S(n86), 
	.B(n2770), 
	.A(n2767));
   MUX2X1 U2462 (.Y(n252), 
	.S(n2989), 
	.B(n2984), 
	.A(n2558));
   XOR2X1 U2463 (.Y(n251), 
	.B(n2988), 
	.A(n2987));
   XOR2X1 U2464 (.Y(n2988), 
	.B(n236), 
	.A(n2823));
   XOR2X1 U2465 (.Y(n250), 
	.B(n233), 
	.A(n235));
   XOR2X1 U2466 (.Y(n236), 
	.B(n2815), 
	.A(n2818));
   AOI21X1 U2467 (.Y(n2990), 
	.C(n2992), 
	.B(DIN[7]), 
	.A(n2991));
   XOR2X1 U2468 (.Y(n235), 
	.B(n2991), 
	.A(DIN[7]));
   XOR2X1 U2469 (.Y(n2991), 
	.B(n238), 
	.A(DIN[4]));
   AOI21X1 U2470 (.Y(n2993), 
	.C(n2995), 
	.B(DIN[3]), 
	.A(n2994));
   XOR2X1 U2471 (.Y(n238), 
	.B(n2994), 
	.A(DIN[3]));
   XOR2X1 U2472 (.Y(n2994), 
	.B(DIN[5]), 
	.A(DIN[6]));
   AOI21X1 U2473 (.Y(n2996), 
	.C(n2998), 
	.B(DIN[0]), 
	.A(n2997));
   XOR2X1 U2474 (.Y(n233), 
	.B(n2997), 
	.A(DIN[0]));
   XOR2X1 U2475 (.Y(n2997), 
	.B(DIN[2]), 
	.A(DIN[1]));
endmodule

